magic
tech sky130B
magscale 1 2
timestamp 1651947127
<< error_p >>
rect -6958 3731 -6898 3850
rect -6878 3731 -6818 3850
rect -7082 2769 -6818 3731
rect -6958 2650 -6898 2769
rect -6878 2650 -6818 2769
rect -6762 2766 -6556 3734
rect -5236 3731 -5176 3850
rect -5156 3731 -5096 3850
rect -5360 2769 -5096 3731
rect -5236 2650 -5176 2769
rect -5156 2650 -5096 2769
rect -5040 2766 -4834 3734
rect -3514 3731 -3454 3850
rect -3434 3731 -3374 3850
rect -3638 2769 -3374 3731
rect -3514 2650 -3454 2769
rect -3434 2650 -3374 2769
rect -3318 2766 -3112 3734
rect -1792 3731 -1732 3850
rect -1712 3731 -1652 3850
rect -1916 2769 -1652 3731
rect -1792 2650 -1732 2769
rect -1712 2650 -1652 2769
rect -1596 2766 -1390 3734
rect -70 3731 -10 3850
rect 10 3731 70 3850
rect -194 2769 70 3731
rect -70 2650 -10 2769
rect 10 2650 70 2769
rect 126 2766 332 3734
rect 1652 3731 1712 3850
rect 1732 3731 1792 3850
rect 1528 2769 1792 3731
rect 1652 2650 1712 2769
rect 1732 2650 1792 2769
rect 1848 2766 2054 3734
rect 3374 3731 3434 3850
rect 3454 3731 3514 3850
rect 3250 2769 3514 3731
rect 3374 2650 3434 2769
rect 3454 2650 3514 2769
rect 3570 2766 3776 3734
rect 5096 3731 5156 3850
rect 5176 3731 5236 3850
rect 4972 2769 5236 3731
rect 5096 2650 5156 2769
rect 5176 2650 5236 2769
rect 5292 2766 5498 3734
rect 6818 3731 6878 3850
rect 6898 3731 6958 3850
rect 6694 2769 6958 3731
rect 6818 2650 6878 2769
rect 6898 2650 6958 2769
rect 7014 2766 7220 3734
rect -6958 2431 -6898 2550
rect -6878 2431 -6818 2550
rect -7082 1469 -6818 2431
rect -6958 1350 -6898 1469
rect -6878 1350 -6818 1469
rect -6762 1466 -6556 2434
rect -5236 2431 -5176 2550
rect -5156 2431 -5096 2550
rect -5360 1469 -5096 2431
rect -5236 1350 -5176 1469
rect -5156 1350 -5096 1469
rect -5040 1466 -4834 2434
rect -3514 2431 -3454 2550
rect -3434 2431 -3374 2550
rect -3638 1469 -3374 2431
rect -3514 1350 -3454 1469
rect -3434 1350 -3374 1469
rect -3318 1466 -3112 2434
rect -1792 2431 -1732 2550
rect -1712 2431 -1652 2550
rect -1916 1469 -1652 2431
rect -1792 1350 -1732 1469
rect -1712 1350 -1652 1469
rect -1596 1466 -1390 2434
rect -70 2431 -10 2550
rect 10 2431 70 2550
rect -194 1469 70 2431
rect -70 1350 -10 1469
rect 10 1350 70 1469
rect 126 1466 332 2434
rect 1652 2431 1712 2550
rect 1732 2431 1792 2550
rect 1528 1469 1792 2431
rect 1652 1350 1712 1469
rect 1732 1350 1792 1469
rect 1848 1466 2054 2434
rect 3374 2431 3434 2550
rect 3454 2431 3514 2550
rect 3250 1469 3514 2431
rect 3374 1350 3434 1469
rect 3454 1350 3514 1469
rect 3570 1466 3776 2434
rect 5096 2431 5156 2550
rect 5176 2431 5236 2550
rect 4972 1469 5236 2431
rect 5096 1350 5156 1469
rect 5176 1350 5236 1469
rect 5292 1466 5498 2434
rect 6818 2431 6878 2550
rect 6898 2431 6958 2550
rect 6694 1469 6958 2431
rect 6818 1350 6878 1469
rect 6898 1350 6958 1469
rect 7014 1466 7220 2434
rect -6958 1131 -6898 1250
rect -6878 1131 -6818 1250
rect -7082 169 -6818 1131
rect -6958 50 -6898 169
rect -6878 50 -6818 169
rect -6762 166 -6556 1134
rect -5236 1131 -5176 1250
rect -5156 1131 -5096 1250
rect -5360 169 -5096 1131
rect -5236 50 -5176 169
rect -5156 50 -5096 169
rect -5040 166 -4834 1134
rect -3514 1131 -3454 1250
rect -3434 1131 -3374 1250
rect -3638 169 -3374 1131
rect -3514 50 -3454 169
rect -3434 50 -3374 169
rect -3318 166 -3112 1134
rect -1792 1131 -1732 1250
rect -1712 1131 -1652 1250
rect -1916 169 -1652 1131
rect -1792 50 -1732 169
rect -1712 50 -1652 169
rect -1596 166 -1390 1134
rect -70 1131 -10 1250
rect 10 1131 70 1250
rect -194 169 70 1131
rect -70 50 -10 169
rect 10 50 70 169
rect 126 166 332 1134
rect 1652 1131 1712 1250
rect 1732 1131 1792 1250
rect 1528 169 1792 1131
rect 1652 50 1712 169
rect 1732 50 1792 169
rect 1848 166 2054 1134
rect 3374 1131 3434 1250
rect 3454 1131 3514 1250
rect 3250 169 3514 1131
rect 3374 50 3434 169
rect 3454 50 3514 169
rect 3570 166 3776 1134
rect 5096 1131 5156 1250
rect 5176 1131 5236 1250
rect 4972 169 5236 1131
rect 5096 50 5156 169
rect 5176 50 5236 169
rect 5292 166 5498 1134
rect 6818 1131 6878 1250
rect 6898 1131 6958 1250
rect 6694 169 6958 1131
rect 6818 50 6878 169
rect 6898 50 6958 169
rect 7014 166 7220 1134
rect -6958 -169 -6898 -50
rect -6878 -169 -6818 -50
rect -7082 -1131 -6818 -169
rect -6958 -1250 -6898 -1131
rect -6878 -1250 -6818 -1131
rect -6762 -1134 -6556 -166
rect -5236 -169 -5176 -50
rect -5156 -169 -5096 -50
rect -5360 -1131 -5096 -169
rect -5236 -1250 -5176 -1131
rect -5156 -1250 -5096 -1131
rect -5040 -1134 -4834 -166
rect -3514 -169 -3454 -50
rect -3434 -169 -3374 -50
rect -3638 -1131 -3374 -169
rect -3514 -1250 -3454 -1131
rect -3434 -1250 -3374 -1131
rect -3318 -1134 -3112 -166
rect -1792 -169 -1732 -50
rect -1712 -169 -1652 -50
rect -1916 -1131 -1652 -169
rect -1792 -1250 -1732 -1131
rect -1712 -1250 -1652 -1131
rect -1596 -1134 -1390 -166
rect -70 -169 -10 -50
rect 10 -169 70 -50
rect -194 -1131 70 -169
rect -70 -1250 -10 -1131
rect 10 -1250 70 -1131
rect 126 -1134 332 -166
rect 1652 -169 1712 -50
rect 1732 -169 1792 -50
rect 1528 -1131 1792 -169
rect 1652 -1250 1712 -1131
rect 1732 -1250 1792 -1131
rect 1848 -1134 2054 -166
rect 3374 -169 3434 -50
rect 3454 -169 3514 -50
rect 3250 -1131 3514 -169
rect 3374 -1250 3434 -1131
rect 3454 -1250 3514 -1131
rect 3570 -1134 3776 -166
rect 5096 -169 5156 -50
rect 5176 -169 5236 -50
rect 4972 -1131 5236 -169
rect 5096 -1250 5156 -1131
rect 5176 -1250 5236 -1131
rect 5292 -1134 5498 -166
rect 6818 -169 6878 -50
rect 6898 -169 6958 -50
rect 6694 -1131 6958 -169
rect 6818 -1250 6878 -1131
rect 6898 -1250 6958 -1131
rect 7014 -1134 7220 -166
rect -6958 -1469 -6898 -1350
rect -6878 -1469 -6818 -1350
rect -7082 -2431 -6818 -1469
rect -6958 -2550 -6898 -2431
rect -6878 -2550 -6818 -2431
rect -6762 -2434 -6556 -1466
rect -5236 -1469 -5176 -1350
rect -5156 -1469 -5096 -1350
rect -5360 -2431 -5096 -1469
rect -5236 -2550 -5176 -2431
rect -5156 -2550 -5096 -2431
rect -5040 -2434 -4834 -1466
rect -3514 -1469 -3454 -1350
rect -3434 -1469 -3374 -1350
rect -3638 -2431 -3374 -1469
rect -3514 -2550 -3454 -2431
rect -3434 -2550 -3374 -2431
rect -3318 -2434 -3112 -1466
rect -1792 -1469 -1732 -1350
rect -1712 -1469 -1652 -1350
rect -1916 -2431 -1652 -1469
rect -1792 -2550 -1732 -2431
rect -1712 -2550 -1652 -2431
rect -1596 -2434 -1390 -1466
rect -70 -1469 -10 -1350
rect 10 -1469 70 -1350
rect -194 -2431 70 -1469
rect -70 -2550 -10 -2431
rect 10 -2550 70 -2431
rect 126 -2434 332 -1466
rect 1652 -1469 1712 -1350
rect 1732 -1469 1792 -1350
rect 1528 -2431 1792 -1469
rect 1652 -2550 1712 -2431
rect 1732 -2550 1792 -2431
rect 1848 -2434 2054 -1466
rect 3374 -1469 3434 -1350
rect 3454 -1469 3514 -1350
rect 3250 -2431 3514 -1469
rect 3374 -2550 3434 -2431
rect 3454 -2550 3514 -2431
rect 3570 -2434 3776 -1466
rect 5096 -1469 5156 -1350
rect 5176 -1469 5236 -1350
rect 4972 -2431 5236 -1469
rect 5096 -2550 5156 -2431
rect 5176 -2550 5236 -2431
rect 5292 -2434 5498 -1466
rect 6818 -1469 6878 -1350
rect 6898 -1469 6958 -1350
rect 6694 -2431 6958 -1469
rect 6818 -2550 6878 -2431
rect 6898 -2550 6958 -2431
rect 7014 -2434 7220 -1466
rect -6958 -2769 -6898 -2650
rect -6878 -2769 -6818 -2650
rect -7082 -3731 -6818 -2769
rect -6958 -3850 -6898 -3731
rect -6878 -3850 -6818 -3731
rect -6762 -3734 -6556 -2766
rect -5236 -2769 -5176 -2650
rect -5156 -2769 -5096 -2650
rect -5360 -3731 -5096 -2769
rect -5236 -3850 -5176 -3731
rect -5156 -3850 -5096 -3731
rect -5040 -3734 -4834 -2766
rect -3514 -2769 -3454 -2650
rect -3434 -2769 -3374 -2650
rect -3638 -3731 -3374 -2769
rect -3514 -3850 -3454 -3731
rect -3434 -3850 -3374 -3731
rect -3318 -3734 -3112 -2766
rect -1792 -2769 -1732 -2650
rect -1712 -2769 -1652 -2650
rect -1916 -3731 -1652 -2769
rect -1792 -3850 -1732 -3731
rect -1712 -3850 -1652 -3731
rect -1596 -3734 -1390 -2766
rect -70 -2769 -10 -2650
rect 10 -2769 70 -2650
rect -194 -3731 70 -2769
rect -70 -3850 -10 -3731
rect 10 -3850 70 -3731
rect 126 -3734 332 -2766
rect 1652 -2769 1712 -2650
rect 1732 -2769 1792 -2650
rect 1528 -3731 1792 -2769
rect 1652 -3850 1712 -3731
rect 1732 -3850 1792 -3731
rect 1848 -3734 2054 -2766
rect 3374 -2769 3434 -2650
rect 3454 -2769 3514 -2650
rect 3250 -3731 3514 -2769
rect 3374 -3850 3434 -3731
rect 3454 -3850 3514 -3731
rect 3570 -3734 3776 -2766
rect 5096 -2769 5156 -2650
rect 5176 -2769 5236 -2650
rect 4972 -3731 5236 -2769
rect 5096 -3850 5156 -3731
rect 5176 -3850 5236 -3731
rect 5292 -3734 5498 -2766
rect 6818 -2769 6878 -2650
rect 6898 -2769 6958 -2650
rect 6694 -3731 6958 -2769
rect 6818 -3850 6878 -3731
rect 6898 -3850 6958 -3731
rect 7014 -3734 7220 -2766
<< metal4 >>
rect -8600 3689 -6898 3850
rect -8600 2811 -7154 3689
rect -6918 2811 -6898 3689
rect -8600 2650 -6898 2811
rect -6878 3689 -5176 3850
rect -6878 2811 -5432 3689
rect -5196 2811 -5176 3689
rect -6878 2650 -5176 2811
rect -5156 3689 -3454 3850
rect -5156 2811 -3710 3689
rect -3474 2811 -3454 3689
rect -5156 2650 -3454 2811
rect -3434 3689 -1732 3850
rect -3434 2811 -1988 3689
rect -1752 2811 -1732 3689
rect -3434 2650 -1732 2811
rect -1712 3689 -10 3850
rect -1712 2811 -266 3689
rect -30 2811 -10 3689
rect -1712 2650 -10 2811
rect 10 3689 1712 3850
rect 10 2811 1456 3689
rect 1692 2811 1712 3689
rect 10 2650 1712 2811
rect 1732 3689 3434 3850
rect 1732 2811 3178 3689
rect 3414 2811 3434 3689
rect 1732 2650 3434 2811
rect 3454 3689 5156 3850
rect 3454 2811 4900 3689
rect 5136 2811 5156 3689
rect 3454 2650 5156 2811
rect 5176 3689 6878 3850
rect 5176 2811 6622 3689
rect 6858 2811 6878 3689
rect 5176 2650 6878 2811
rect 6898 3689 8600 3850
rect 6898 2811 8344 3689
rect 8580 2811 8600 3689
rect 6898 2650 8600 2811
rect -8600 2389 -6898 2550
rect -8600 1511 -7154 2389
rect -6918 1511 -6898 2389
rect -8600 1350 -6898 1511
rect -6878 2389 -5176 2550
rect -6878 1511 -5432 2389
rect -5196 1511 -5176 2389
rect -6878 1350 -5176 1511
rect -5156 2389 -3454 2550
rect -5156 1511 -3710 2389
rect -3474 1511 -3454 2389
rect -5156 1350 -3454 1511
rect -3434 2389 -1732 2550
rect -3434 1511 -1988 2389
rect -1752 1511 -1732 2389
rect -3434 1350 -1732 1511
rect -1712 2389 -10 2550
rect -1712 1511 -266 2389
rect -30 1511 -10 2389
rect -1712 1350 -10 1511
rect 10 2389 1712 2550
rect 10 1511 1456 2389
rect 1692 1511 1712 2389
rect 10 1350 1712 1511
rect 1732 2389 3434 2550
rect 1732 1511 3178 2389
rect 3414 1511 3434 2389
rect 1732 1350 3434 1511
rect 3454 2389 5156 2550
rect 3454 1511 4900 2389
rect 5136 1511 5156 2389
rect 3454 1350 5156 1511
rect 5176 2389 6878 2550
rect 5176 1511 6622 2389
rect 6858 1511 6878 2389
rect 5176 1350 6878 1511
rect 6898 2389 8600 2550
rect 6898 1511 8344 2389
rect 8580 1511 8600 2389
rect 6898 1350 8600 1511
rect -8600 1089 -6898 1250
rect -8600 211 -7154 1089
rect -6918 211 -6898 1089
rect -8600 50 -6898 211
rect -6878 1089 -5176 1250
rect -6878 211 -5432 1089
rect -5196 211 -5176 1089
rect -6878 50 -5176 211
rect -5156 1089 -3454 1250
rect -5156 211 -3710 1089
rect -3474 211 -3454 1089
rect -5156 50 -3454 211
rect -3434 1089 -1732 1250
rect -3434 211 -1988 1089
rect -1752 211 -1732 1089
rect -3434 50 -1732 211
rect -1712 1089 -10 1250
rect -1712 211 -266 1089
rect -30 211 -10 1089
rect -1712 50 -10 211
rect 10 1089 1712 1250
rect 10 211 1456 1089
rect 1692 211 1712 1089
rect 10 50 1712 211
rect 1732 1089 3434 1250
rect 1732 211 3178 1089
rect 3414 211 3434 1089
rect 1732 50 3434 211
rect 3454 1089 5156 1250
rect 3454 211 4900 1089
rect 5136 211 5156 1089
rect 3454 50 5156 211
rect 5176 1089 6878 1250
rect 5176 211 6622 1089
rect 6858 211 6878 1089
rect 5176 50 6878 211
rect 6898 1089 8600 1250
rect 6898 211 8344 1089
rect 8580 211 8600 1089
rect 6898 50 8600 211
rect -8600 -211 -6898 -50
rect -8600 -1089 -7154 -211
rect -6918 -1089 -6898 -211
rect -8600 -1250 -6898 -1089
rect -6878 -211 -5176 -50
rect -6878 -1089 -5432 -211
rect -5196 -1089 -5176 -211
rect -6878 -1250 -5176 -1089
rect -5156 -211 -3454 -50
rect -5156 -1089 -3710 -211
rect -3474 -1089 -3454 -211
rect -5156 -1250 -3454 -1089
rect -3434 -211 -1732 -50
rect -3434 -1089 -1988 -211
rect -1752 -1089 -1732 -211
rect -3434 -1250 -1732 -1089
rect -1712 -211 -10 -50
rect -1712 -1089 -266 -211
rect -30 -1089 -10 -211
rect -1712 -1250 -10 -1089
rect 10 -211 1712 -50
rect 10 -1089 1456 -211
rect 1692 -1089 1712 -211
rect 10 -1250 1712 -1089
rect 1732 -211 3434 -50
rect 1732 -1089 3178 -211
rect 3414 -1089 3434 -211
rect 1732 -1250 3434 -1089
rect 3454 -211 5156 -50
rect 3454 -1089 4900 -211
rect 5136 -1089 5156 -211
rect 3454 -1250 5156 -1089
rect 5176 -211 6878 -50
rect 5176 -1089 6622 -211
rect 6858 -1089 6878 -211
rect 5176 -1250 6878 -1089
rect 6898 -211 8600 -50
rect 6898 -1089 8344 -211
rect 8580 -1089 8600 -211
rect 6898 -1250 8600 -1089
rect -8600 -1511 -6898 -1350
rect -8600 -2389 -7154 -1511
rect -6918 -2389 -6898 -1511
rect -8600 -2550 -6898 -2389
rect -6878 -1511 -5176 -1350
rect -6878 -2389 -5432 -1511
rect -5196 -2389 -5176 -1511
rect -6878 -2550 -5176 -2389
rect -5156 -1511 -3454 -1350
rect -5156 -2389 -3710 -1511
rect -3474 -2389 -3454 -1511
rect -5156 -2550 -3454 -2389
rect -3434 -1511 -1732 -1350
rect -3434 -2389 -1988 -1511
rect -1752 -2389 -1732 -1511
rect -3434 -2550 -1732 -2389
rect -1712 -1511 -10 -1350
rect -1712 -2389 -266 -1511
rect -30 -2389 -10 -1511
rect -1712 -2550 -10 -2389
rect 10 -1511 1712 -1350
rect 10 -2389 1456 -1511
rect 1692 -2389 1712 -1511
rect 10 -2550 1712 -2389
rect 1732 -1511 3434 -1350
rect 1732 -2389 3178 -1511
rect 3414 -2389 3434 -1511
rect 1732 -2550 3434 -2389
rect 3454 -1511 5156 -1350
rect 3454 -2389 4900 -1511
rect 5136 -2389 5156 -1511
rect 3454 -2550 5156 -2389
rect 5176 -1511 6878 -1350
rect 5176 -2389 6622 -1511
rect 6858 -2389 6878 -1511
rect 5176 -2550 6878 -2389
rect 6898 -1511 8600 -1350
rect 6898 -2389 8344 -1511
rect 8580 -2389 8600 -1511
rect 6898 -2550 8600 -2389
rect -8600 -2811 -6898 -2650
rect -8600 -3689 -7154 -2811
rect -6918 -3689 -6898 -2811
rect -8600 -3850 -6898 -3689
rect -6878 -2811 -5176 -2650
rect -6878 -3689 -5432 -2811
rect -5196 -3689 -5176 -2811
rect -6878 -3850 -5176 -3689
rect -5156 -2811 -3454 -2650
rect -5156 -3689 -3710 -2811
rect -3474 -3689 -3454 -2811
rect -5156 -3850 -3454 -3689
rect -3434 -2811 -1732 -2650
rect -3434 -3689 -1988 -2811
rect -1752 -3689 -1732 -2811
rect -3434 -3850 -1732 -3689
rect -1712 -2811 -10 -2650
rect -1712 -3689 -266 -2811
rect -30 -3689 -10 -2811
rect -1712 -3850 -10 -3689
rect 10 -2811 1712 -2650
rect 10 -3689 1456 -2811
rect 1692 -3689 1712 -2811
rect 10 -3850 1712 -3689
rect 1732 -2811 3434 -2650
rect 1732 -3689 3178 -2811
rect 3414 -3689 3434 -2811
rect 1732 -3850 3434 -3689
rect 3454 -2811 5156 -2650
rect 3454 -3689 4900 -2811
rect 5136 -3689 5156 -2811
rect 3454 -3850 5156 -3689
rect 5176 -2811 6878 -2650
rect 5176 -3689 6622 -2811
rect 6858 -3689 6878 -2811
rect 5176 -3850 6878 -3689
rect 6898 -2811 8600 -2650
rect 6898 -3689 8344 -2811
rect 8580 -3689 8600 -2811
rect 6898 -3850 8600 -3689
<< via4 >>
rect -7154 2811 -6918 3689
rect -5432 2811 -5196 3689
rect -3710 2811 -3474 3689
rect -1988 2811 -1752 3689
rect -266 2811 -30 3689
rect 1456 2811 1692 3689
rect 3178 2811 3414 3689
rect 4900 2811 5136 3689
rect 6622 2811 6858 3689
rect 8344 2811 8580 3689
rect -7154 1511 -6918 2389
rect -5432 1511 -5196 2389
rect -3710 1511 -3474 2389
rect -1988 1511 -1752 2389
rect -266 1511 -30 2389
rect 1456 1511 1692 2389
rect 3178 1511 3414 2389
rect 4900 1511 5136 2389
rect 6622 1511 6858 2389
rect 8344 1511 8580 2389
rect -7154 211 -6918 1089
rect -5432 211 -5196 1089
rect -3710 211 -3474 1089
rect -1988 211 -1752 1089
rect -266 211 -30 1089
rect 1456 211 1692 1089
rect 3178 211 3414 1089
rect 4900 211 5136 1089
rect 6622 211 6858 1089
rect 8344 211 8580 1089
rect -7154 -1089 -6918 -211
rect -5432 -1089 -5196 -211
rect -3710 -1089 -3474 -211
rect -1988 -1089 -1752 -211
rect -266 -1089 -30 -211
rect 1456 -1089 1692 -211
rect 3178 -1089 3414 -211
rect 4900 -1089 5136 -211
rect 6622 -1089 6858 -211
rect 8344 -1089 8580 -211
rect -7154 -2389 -6918 -1511
rect -5432 -2389 -5196 -1511
rect -3710 -2389 -3474 -1511
rect -1988 -2389 -1752 -1511
rect -266 -2389 -30 -1511
rect 1456 -2389 1692 -1511
rect 3178 -2389 3414 -1511
rect 4900 -2389 5136 -1511
rect 6622 -2389 6858 -1511
rect 8344 -2389 8580 -1511
rect -7154 -3689 -6918 -2811
rect -5432 -3689 -5196 -2811
rect -3710 -3689 -3474 -2811
rect -1988 -3689 -1752 -2811
rect -266 -3689 -30 -2811
rect 1456 -3689 1692 -2811
rect 3178 -3689 3414 -2811
rect 4900 -3689 5136 -2811
rect 6622 -3689 6858 -2811
rect 8344 -3689 8580 -2811
<< mimcap2 >>
rect -8500 3710 -7500 3750
rect -8500 2790 -8460 3710
rect -7540 2790 -7500 3710
rect -8500 2750 -7500 2790
rect -6778 3710 -5778 3750
rect -6778 2790 -6738 3710
rect -5818 2790 -5778 3710
rect -6778 2750 -5778 2790
rect -5056 3710 -4056 3750
rect -5056 2790 -5016 3710
rect -4096 2790 -4056 3710
rect -5056 2750 -4056 2790
rect -3334 3710 -2334 3750
rect -3334 2790 -3294 3710
rect -2374 2790 -2334 3710
rect -3334 2750 -2334 2790
rect -1612 3710 -612 3750
rect -1612 2790 -1572 3710
rect -652 2790 -612 3710
rect -1612 2750 -612 2790
rect 110 3710 1110 3750
rect 110 2790 150 3710
rect 1070 2790 1110 3710
rect 110 2750 1110 2790
rect 1832 3710 2832 3750
rect 1832 2790 1872 3710
rect 2792 2790 2832 3710
rect 1832 2750 2832 2790
rect 3554 3710 4554 3750
rect 3554 2790 3594 3710
rect 4514 2790 4554 3710
rect 3554 2750 4554 2790
rect 5276 3710 6276 3750
rect 5276 2790 5316 3710
rect 6236 2790 6276 3710
rect 5276 2750 6276 2790
rect 6998 3710 7998 3750
rect 6998 2790 7038 3710
rect 7958 2790 7998 3710
rect 6998 2750 7998 2790
rect -8500 2410 -7500 2450
rect -8500 1490 -8460 2410
rect -7540 1490 -7500 2410
rect -8500 1450 -7500 1490
rect -6778 2410 -5778 2450
rect -6778 1490 -6738 2410
rect -5818 1490 -5778 2410
rect -6778 1450 -5778 1490
rect -5056 2410 -4056 2450
rect -5056 1490 -5016 2410
rect -4096 1490 -4056 2410
rect -5056 1450 -4056 1490
rect -3334 2410 -2334 2450
rect -3334 1490 -3294 2410
rect -2374 1490 -2334 2410
rect -3334 1450 -2334 1490
rect -1612 2410 -612 2450
rect -1612 1490 -1572 2410
rect -652 1490 -612 2410
rect -1612 1450 -612 1490
rect 110 2410 1110 2450
rect 110 1490 150 2410
rect 1070 1490 1110 2410
rect 110 1450 1110 1490
rect 1832 2410 2832 2450
rect 1832 1490 1872 2410
rect 2792 1490 2832 2410
rect 1832 1450 2832 1490
rect 3554 2410 4554 2450
rect 3554 1490 3594 2410
rect 4514 1490 4554 2410
rect 3554 1450 4554 1490
rect 5276 2410 6276 2450
rect 5276 1490 5316 2410
rect 6236 1490 6276 2410
rect 5276 1450 6276 1490
rect 6998 2410 7998 2450
rect 6998 1490 7038 2410
rect 7958 1490 7998 2410
rect 6998 1450 7998 1490
rect -8500 1110 -7500 1150
rect -8500 190 -8460 1110
rect -7540 190 -7500 1110
rect -8500 150 -7500 190
rect -6778 1110 -5778 1150
rect -6778 190 -6738 1110
rect -5818 190 -5778 1110
rect -6778 150 -5778 190
rect -5056 1110 -4056 1150
rect -5056 190 -5016 1110
rect -4096 190 -4056 1110
rect -5056 150 -4056 190
rect -3334 1110 -2334 1150
rect -3334 190 -3294 1110
rect -2374 190 -2334 1110
rect -3334 150 -2334 190
rect -1612 1110 -612 1150
rect -1612 190 -1572 1110
rect -652 190 -612 1110
rect -1612 150 -612 190
rect 110 1110 1110 1150
rect 110 190 150 1110
rect 1070 190 1110 1110
rect 110 150 1110 190
rect 1832 1110 2832 1150
rect 1832 190 1872 1110
rect 2792 190 2832 1110
rect 1832 150 2832 190
rect 3554 1110 4554 1150
rect 3554 190 3594 1110
rect 4514 190 4554 1110
rect 3554 150 4554 190
rect 5276 1110 6276 1150
rect 5276 190 5316 1110
rect 6236 190 6276 1110
rect 5276 150 6276 190
rect 6998 1110 7998 1150
rect 6998 190 7038 1110
rect 7958 190 7998 1110
rect 6998 150 7998 190
rect -8500 -190 -7500 -150
rect -8500 -1110 -8460 -190
rect -7540 -1110 -7500 -190
rect -8500 -1150 -7500 -1110
rect -6778 -190 -5778 -150
rect -6778 -1110 -6738 -190
rect -5818 -1110 -5778 -190
rect -6778 -1150 -5778 -1110
rect -5056 -190 -4056 -150
rect -5056 -1110 -5016 -190
rect -4096 -1110 -4056 -190
rect -5056 -1150 -4056 -1110
rect -3334 -190 -2334 -150
rect -3334 -1110 -3294 -190
rect -2374 -1110 -2334 -190
rect -3334 -1150 -2334 -1110
rect -1612 -190 -612 -150
rect -1612 -1110 -1572 -190
rect -652 -1110 -612 -190
rect -1612 -1150 -612 -1110
rect 110 -190 1110 -150
rect 110 -1110 150 -190
rect 1070 -1110 1110 -190
rect 110 -1150 1110 -1110
rect 1832 -190 2832 -150
rect 1832 -1110 1872 -190
rect 2792 -1110 2832 -190
rect 1832 -1150 2832 -1110
rect 3554 -190 4554 -150
rect 3554 -1110 3594 -190
rect 4514 -1110 4554 -190
rect 3554 -1150 4554 -1110
rect 5276 -190 6276 -150
rect 5276 -1110 5316 -190
rect 6236 -1110 6276 -190
rect 5276 -1150 6276 -1110
rect 6998 -190 7998 -150
rect 6998 -1110 7038 -190
rect 7958 -1110 7998 -190
rect 6998 -1150 7998 -1110
rect -8500 -1490 -7500 -1450
rect -8500 -2410 -8460 -1490
rect -7540 -2410 -7500 -1490
rect -8500 -2450 -7500 -2410
rect -6778 -1490 -5778 -1450
rect -6778 -2410 -6738 -1490
rect -5818 -2410 -5778 -1490
rect -6778 -2450 -5778 -2410
rect -5056 -1490 -4056 -1450
rect -5056 -2410 -5016 -1490
rect -4096 -2410 -4056 -1490
rect -5056 -2450 -4056 -2410
rect -3334 -1490 -2334 -1450
rect -3334 -2410 -3294 -1490
rect -2374 -2410 -2334 -1490
rect -3334 -2450 -2334 -2410
rect -1612 -1490 -612 -1450
rect -1612 -2410 -1572 -1490
rect -652 -2410 -612 -1490
rect -1612 -2450 -612 -2410
rect 110 -1490 1110 -1450
rect 110 -2410 150 -1490
rect 1070 -2410 1110 -1490
rect 110 -2450 1110 -2410
rect 1832 -1490 2832 -1450
rect 1832 -2410 1872 -1490
rect 2792 -2410 2832 -1490
rect 1832 -2450 2832 -2410
rect 3554 -1490 4554 -1450
rect 3554 -2410 3594 -1490
rect 4514 -2410 4554 -1490
rect 3554 -2450 4554 -2410
rect 5276 -1490 6276 -1450
rect 5276 -2410 5316 -1490
rect 6236 -2410 6276 -1490
rect 5276 -2450 6276 -2410
rect 6998 -1490 7998 -1450
rect 6998 -2410 7038 -1490
rect 7958 -2410 7998 -1490
rect 6998 -2450 7998 -2410
rect -8500 -2790 -7500 -2750
rect -8500 -3710 -8460 -2790
rect -7540 -3710 -7500 -2790
rect -8500 -3750 -7500 -3710
rect -6778 -2790 -5778 -2750
rect -6778 -3710 -6738 -2790
rect -5818 -3710 -5778 -2790
rect -6778 -3750 -5778 -3710
rect -5056 -2790 -4056 -2750
rect -5056 -3710 -5016 -2790
rect -4096 -3710 -4056 -2790
rect -5056 -3750 -4056 -3710
rect -3334 -2790 -2334 -2750
rect -3334 -3710 -3294 -2790
rect -2374 -3710 -2334 -2790
rect -3334 -3750 -2334 -3710
rect -1612 -2790 -612 -2750
rect -1612 -3710 -1572 -2790
rect -652 -3710 -612 -2790
rect -1612 -3750 -612 -3710
rect 110 -2790 1110 -2750
rect 110 -3710 150 -2790
rect 1070 -3710 1110 -2790
rect 110 -3750 1110 -3710
rect 1832 -2790 2832 -2750
rect 1832 -3710 1872 -2790
rect 2792 -3710 2832 -2790
rect 1832 -3750 2832 -3710
rect 3554 -2790 4554 -2750
rect 3554 -3710 3594 -2790
rect 4514 -3710 4554 -2790
rect 3554 -3750 4554 -3710
rect 5276 -2790 6276 -2750
rect 5276 -3710 5316 -2790
rect 6236 -3710 6276 -2790
rect 5276 -3750 6276 -3710
rect 6998 -2790 7998 -2750
rect 6998 -3710 7038 -2790
rect 7958 -3710 7998 -2790
rect 6998 -3750 7998 -3710
<< mimcap2contact >>
rect -8460 2790 -7540 3710
rect -6738 2790 -5818 3710
rect -5016 2790 -4096 3710
rect -3294 2790 -2374 3710
rect -1572 2790 -652 3710
rect 150 2790 1070 3710
rect 1872 2790 2792 3710
rect 3594 2790 4514 3710
rect 5316 2790 6236 3710
rect 7038 2790 7958 3710
rect -8460 1490 -7540 2410
rect -6738 1490 -5818 2410
rect -5016 1490 -4096 2410
rect -3294 1490 -2374 2410
rect -1572 1490 -652 2410
rect 150 1490 1070 2410
rect 1872 1490 2792 2410
rect 3594 1490 4514 2410
rect 5316 1490 6236 2410
rect 7038 1490 7958 2410
rect -8460 190 -7540 1110
rect -6738 190 -5818 1110
rect -5016 190 -4096 1110
rect -3294 190 -2374 1110
rect -1572 190 -652 1110
rect 150 190 1070 1110
rect 1872 190 2792 1110
rect 3594 190 4514 1110
rect 5316 190 6236 1110
rect 7038 190 7958 1110
rect -8460 -1110 -7540 -190
rect -6738 -1110 -5818 -190
rect -5016 -1110 -4096 -190
rect -3294 -1110 -2374 -190
rect -1572 -1110 -652 -190
rect 150 -1110 1070 -190
rect 1872 -1110 2792 -190
rect 3594 -1110 4514 -190
rect 5316 -1110 6236 -190
rect 7038 -1110 7958 -190
rect -8460 -2410 -7540 -1490
rect -6738 -2410 -5818 -1490
rect -5016 -2410 -4096 -1490
rect -3294 -2410 -2374 -1490
rect -1572 -2410 -652 -1490
rect 150 -2410 1070 -1490
rect 1872 -2410 2792 -1490
rect 3594 -2410 4514 -1490
rect 5316 -2410 6236 -1490
rect 7038 -2410 7958 -1490
rect -8460 -3710 -7540 -2790
rect -6738 -3710 -5818 -2790
rect -5016 -3710 -4096 -2790
rect -3294 -3710 -2374 -2790
rect -1572 -3710 -652 -2790
rect 150 -3710 1070 -2790
rect 1872 -3710 2792 -2790
rect 3594 -3710 4514 -2790
rect 5316 -3710 6236 -2790
rect 7038 -3710 7958 -2790
<< metal5 >>
rect -8160 3734 -7840 3900
rect -6438 3734 -6118 3900
rect -4716 3734 -4396 3900
rect -2994 3734 -2674 3900
rect -1272 3734 -952 3900
rect 450 3734 770 3900
rect 2172 3734 2492 3900
rect 3894 3734 4214 3900
rect 5616 3734 5936 3900
rect 7338 3734 7658 3900
rect -8484 3710 -7516 3734
rect -8484 2790 -8460 3710
rect -7540 2790 -7516 3710
rect -8484 2766 -7516 2790
rect -7196 3689 -6876 3731
rect -7196 2811 -7154 3689
rect -6918 2811 -6876 3689
rect -7196 2769 -6876 2811
rect -6762 3710 -5794 3734
rect -6762 2790 -6738 3710
rect -5818 2790 -5794 3710
rect -6762 2766 -5794 2790
rect -5474 3689 -5154 3731
rect -5474 2811 -5432 3689
rect -5196 2811 -5154 3689
rect -5474 2769 -5154 2811
rect -5040 3710 -4072 3734
rect -5040 2790 -5016 3710
rect -4096 2790 -4072 3710
rect -5040 2766 -4072 2790
rect -3752 3689 -3432 3731
rect -3752 2811 -3710 3689
rect -3474 2811 -3432 3689
rect -3752 2769 -3432 2811
rect -3318 3710 -2350 3734
rect -3318 2790 -3294 3710
rect -2374 2790 -2350 3710
rect -3318 2766 -2350 2790
rect -2030 3689 -1710 3731
rect -2030 2811 -1988 3689
rect -1752 2811 -1710 3689
rect -2030 2769 -1710 2811
rect -1596 3710 -628 3734
rect -1596 2790 -1572 3710
rect -652 2790 -628 3710
rect -1596 2766 -628 2790
rect -308 3689 12 3731
rect -308 2811 -266 3689
rect -30 2811 12 3689
rect -308 2769 12 2811
rect 126 3710 1094 3734
rect 126 2790 150 3710
rect 1070 2790 1094 3710
rect 126 2766 1094 2790
rect 1414 3689 1734 3731
rect 1414 2811 1456 3689
rect 1692 2811 1734 3689
rect 1414 2769 1734 2811
rect 1848 3710 2816 3734
rect 1848 2790 1872 3710
rect 2792 2790 2816 3710
rect 1848 2766 2816 2790
rect 3136 3689 3456 3731
rect 3136 2811 3178 3689
rect 3414 2811 3456 3689
rect 3136 2769 3456 2811
rect 3570 3710 4538 3734
rect 3570 2790 3594 3710
rect 4514 2790 4538 3710
rect 3570 2766 4538 2790
rect 4858 3689 5178 3731
rect 4858 2811 4900 3689
rect 5136 2811 5178 3689
rect 4858 2769 5178 2811
rect 5292 3710 6260 3734
rect 5292 2790 5316 3710
rect 6236 2790 6260 3710
rect 5292 2766 6260 2790
rect 6580 3689 6900 3731
rect 6580 2811 6622 3689
rect 6858 2811 6900 3689
rect 6580 2769 6900 2811
rect 7014 3710 7982 3734
rect 7014 2790 7038 3710
rect 7958 2790 7982 3710
rect 7014 2766 7982 2790
rect 8302 3689 8622 3731
rect 8302 2811 8344 3689
rect 8580 2811 8622 3689
rect 8302 2769 8622 2811
rect -8160 2434 -7840 2766
rect -6438 2434 -6118 2766
rect -4716 2434 -4396 2766
rect -2994 2434 -2674 2766
rect -1272 2434 -952 2766
rect 450 2434 770 2766
rect 2172 2434 2492 2766
rect 3894 2434 4214 2766
rect 5616 2434 5936 2766
rect 7338 2434 7658 2766
rect -8484 2410 -7516 2434
rect -8484 1490 -8460 2410
rect -7540 1490 -7516 2410
rect -8484 1466 -7516 1490
rect -7196 2389 -6876 2431
rect -7196 1511 -7154 2389
rect -6918 1511 -6876 2389
rect -7196 1469 -6876 1511
rect -6762 2410 -5794 2434
rect -6762 1490 -6738 2410
rect -5818 1490 -5794 2410
rect -6762 1466 -5794 1490
rect -5474 2389 -5154 2431
rect -5474 1511 -5432 2389
rect -5196 1511 -5154 2389
rect -5474 1469 -5154 1511
rect -5040 2410 -4072 2434
rect -5040 1490 -5016 2410
rect -4096 1490 -4072 2410
rect -5040 1466 -4072 1490
rect -3752 2389 -3432 2431
rect -3752 1511 -3710 2389
rect -3474 1511 -3432 2389
rect -3752 1469 -3432 1511
rect -3318 2410 -2350 2434
rect -3318 1490 -3294 2410
rect -2374 1490 -2350 2410
rect -3318 1466 -2350 1490
rect -2030 2389 -1710 2431
rect -2030 1511 -1988 2389
rect -1752 1511 -1710 2389
rect -2030 1469 -1710 1511
rect -1596 2410 -628 2434
rect -1596 1490 -1572 2410
rect -652 1490 -628 2410
rect -1596 1466 -628 1490
rect -308 2389 12 2431
rect -308 1511 -266 2389
rect -30 1511 12 2389
rect -308 1469 12 1511
rect 126 2410 1094 2434
rect 126 1490 150 2410
rect 1070 1490 1094 2410
rect 126 1466 1094 1490
rect 1414 2389 1734 2431
rect 1414 1511 1456 2389
rect 1692 1511 1734 2389
rect 1414 1469 1734 1511
rect 1848 2410 2816 2434
rect 1848 1490 1872 2410
rect 2792 1490 2816 2410
rect 1848 1466 2816 1490
rect 3136 2389 3456 2431
rect 3136 1511 3178 2389
rect 3414 1511 3456 2389
rect 3136 1469 3456 1511
rect 3570 2410 4538 2434
rect 3570 1490 3594 2410
rect 4514 1490 4538 2410
rect 3570 1466 4538 1490
rect 4858 2389 5178 2431
rect 4858 1511 4900 2389
rect 5136 1511 5178 2389
rect 4858 1469 5178 1511
rect 5292 2410 6260 2434
rect 5292 1490 5316 2410
rect 6236 1490 6260 2410
rect 5292 1466 6260 1490
rect 6580 2389 6900 2431
rect 6580 1511 6622 2389
rect 6858 1511 6900 2389
rect 6580 1469 6900 1511
rect 7014 2410 7982 2434
rect 7014 1490 7038 2410
rect 7958 1490 7982 2410
rect 7014 1466 7982 1490
rect 8302 2389 8622 2431
rect 8302 1511 8344 2389
rect 8580 1511 8622 2389
rect 8302 1469 8622 1511
rect -8160 1134 -7840 1466
rect -6438 1134 -6118 1466
rect -4716 1134 -4396 1466
rect -2994 1134 -2674 1466
rect -1272 1134 -952 1466
rect 450 1134 770 1466
rect 2172 1134 2492 1466
rect 3894 1134 4214 1466
rect 5616 1134 5936 1466
rect 7338 1134 7658 1466
rect -8484 1110 -7516 1134
rect -8484 190 -8460 1110
rect -7540 190 -7516 1110
rect -8484 166 -7516 190
rect -7196 1089 -6876 1131
rect -7196 211 -7154 1089
rect -6918 211 -6876 1089
rect -7196 169 -6876 211
rect -6762 1110 -5794 1134
rect -6762 190 -6738 1110
rect -5818 190 -5794 1110
rect -6762 166 -5794 190
rect -5474 1089 -5154 1131
rect -5474 211 -5432 1089
rect -5196 211 -5154 1089
rect -5474 169 -5154 211
rect -5040 1110 -4072 1134
rect -5040 190 -5016 1110
rect -4096 190 -4072 1110
rect -5040 166 -4072 190
rect -3752 1089 -3432 1131
rect -3752 211 -3710 1089
rect -3474 211 -3432 1089
rect -3752 169 -3432 211
rect -3318 1110 -2350 1134
rect -3318 190 -3294 1110
rect -2374 190 -2350 1110
rect -3318 166 -2350 190
rect -2030 1089 -1710 1131
rect -2030 211 -1988 1089
rect -1752 211 -1710 1089
rect -2030 169 -1710 211
rect -1596 1110 -628 1134
rect -1596 190 -1572 1110
rect -652 190 -628 1110
rect -1596 166 -628 190
rect -308 1089 12 1131
rect -308 211 -266 1089
rect -30 211 12 1089
rect -308 169 12 211
rect 126 1110 1094 1134
rect 126 190 150 1110
rect 1070 190 1094 1110
rect 126 166 1094 190
rect 1414 1089 1734 1131
rect 1414 211 1456 1089
rect 1692 211 1734 1089
rect 1414 169 1734 211
rect 1848 1110 2816 1134
rect 1848 190 1872 1110
rect 2792 190 2816 1110
rect 1848 166 2816 190
rect 3136 1089 3456 1131
rect 3136 211 3178 1089
rect 3414 211 3456 1089
rect 3136 169 3456 211
rect 3570 1110 4538 1134
rect 3570 190 3594 1110
rect 4514 190 4538 1110
rect 3570 166 4538 190
rect 4858 1089 5178 1131
rect 4858 211 4900 1089
rect 5136 211 5178 1089
rect 4858 169 5178 211
rect 5292 1110 6260 1134
rect 5292 190 5316 1110
rect 6236 190 6260 1110
rect 5292 166 6260 190
rect 6580 1089 6900 1131
rect 6580 211 6622 1089
rect 6858 211 6900 1089
rect 6580 169 6900 211
rect 7014 1110 7982 1134
rect 7014 190 7038 1110
rect 7958 190 7982 1110
rect 7014 166 7982 190
rect 8302 1089 8622 1131
rect 8302 211 8344 1089
rect 8580 211 8622 1089
rect 8302 169 8622 211
rect -8160 -166 -7840 166
rect -6438 -166 -6118 166
rect -4716 -166 -4396 166
rect -2994 -166 -2674 166
rect -1272 -166 -952 166
rect 450 -166 770 166
rect 2172 -166 2492 166
rect 3894 -166 4214 166
rect 5616 -166 5936 166
rect 7338 -166 7658 166
rect -8484 -190 -7516 -166
rect -8484 -1110 -8460 -190
rect -7540 -1110 -7516 -190
rect -8484 -1134 -7516 -1110
rect -7196 -211 -6876 -169
rect -7196 -1089 -7154 -211
rect -6918 -1089 -6876 -211
rect -7196 -1131 -6876 -1089
rect -6762 -190 -5794 -166
rect -6762 -1110 -6738 -190
rect -5818 -1110 -5794 -190
rect -6762 -1134 -5794 -1110
rect -5474 -211 -5154 -169
rect -5474 -1089 -5432 -211
rect -5196 -1089 -5154 -211
rect -5474 -1131 -5154 -1089
rect -5040 -190 -4072 -166
rect -5040 -1110 -5016 -190
rect -4096 -1110 -4072 -190
rect -5040 -1134 -4072 -1110
rect -3752 -211 -3432 -169
rect -3752 -1089 -3710 -211
rect -3474 -1089 -3432 -211
rect -3752 -1131 -3432 -1089
rect -3318 -190 -2350 -166
rect -3318 -1110 -3294 -190
rect -2374 -1110 -2350 -190
rect -3318 -1134 -2350 -1110
rect -2030 -211 -1710 -169
rect -2030 -1089 -1988 -211
rect -1752 -1089 -1710 -211
rect -2030 -1131 -1710 -1089
rect -1596 -190 -628 -166
rect -1596 -1110 -1572 -190
rect -652 -1110 -628 -190
rect -1596 -1134 -628 -1110
rect -308 -211 12 -169
rect -308 -1089 -266 -211
rect -30 -1089 12 -211
rect -308 -1131 12 -1089
rect 126 -190 1094 -166
rect 126 -1110 150 -190
rect 1070 -1110 1094 -190
rect 126 -1134 1094 -1110
rect 1414 -211 1734 -169
rect 1414 -1089 1456 -211
rect 1692 -1089 1734 -211
rect 1414 -1131 1734 -1089
rect 1848 -190 2816 -166
rect 1848 -1110 1872 -190
rect 2792 -1110 2816 -190
rect 1848 -1134 2816 -1110
rect 3136 -211 3456 -169
rect 3136 -1089 3178 -211
rect 3414 -1089 3456 -211
rect 3136 -1131 3456 -1089
rect 3570 -190 4538 -166
rect 3570 -1110 3594 -190
rect 4514 -1110 4538 -190
rect 3570 -1134 4538 -1110
rect 4858 -211 5178 -169
rect 4858 -1089 4900 -211
rect 5136 -1089 5178 -211
rect 4858 -1131 5178 -1089
rect 5292 -190 6260 -166
rect 5292 -1110 5316 -190
rect 6236 -1110 6260 -190
rect 5292 -1134 6260 -1110
rect 6580 -211 6900 -169
rect 6580 -1089 6622 -211
rect 6858 -1089 6900 -211
rect 6580 -1131 6900 -1089
rect 7014 -190 7982 -166
rect 7014 -1110 7038 -190
rect 7958 -1110 7982 -190
rect 7014 -1134 7982 -1110
rect 8302 -211 8622 -169
rect 8302 -1089 8344 -211
rect 8580 -1089 8622 -211
rect 8302 -1131 8622 -1089
rect -8160 -1466 -7840 -1134
rect -6438 -1466 -6118 -1134
rect -4716 -1466 -4396 -1134
rect -2994 -1466 -2674 -1134
rect -1272 -1466 -952 -1134
rect 450 -1466 770 -1134
rect 2172 -1466 2492 -1134
rect 3894 -1466 4214 -1134
rect 5616 -1466 5936 -1134
rect 7338 -1466 7658 -1134
rect -8484 -1490 -7516 -1466
rect -8484 -2410 -8460 -1490
rect -7540 -2410 -7516 -1490
rect -8484 -2434 -7516 -2410
rect -7196 -1511 -6876 -1469
rect -7196 -2389 -7154 -1511
rect -6918 -2389 -6876 -1511
rect -7196 -2431 -6876 -2389
rect -6762 -1490 -5794 -1466
rect -6762 -2410 -6738 -1490
rect -5818 -2410 -5794 -1490
rect -6762 -2434 -5794 -2410
rect -5474 -1511 -5154 -1469
rect -5474 -2389 -5432 -1511
rect -5196 -2389 -5154 -1511
rect -5474 -2431 -5154 -2389
rect -5040 -1490 -4072 -1466
rect -5040 -2410 -5016 -1490
rect -4096 -2410 -4072 -1490
rect -5040 -2434 -4072 -2410
rect -3752 -1511 -3432 -1469
rect -3752 -2389 -3710 -1511
rect -3474 -2389 -3432 -1511
rect -3752 -2431 -3432 -2389
rect -3318 -1490 -2350 -1466
rect -3318 -2410 -3294 -1490
rect -2374 -2410 -2350 -1490
rect -3318 -2434 -2350 -2410
rect -2030 -1511 -1710 -1469
rect -2030 -2389 -1988 -1511
rect -1752 -2389 -1710 -1511
rect -2030 -2431 -1710 -2389
rect -1596 -1490 -628 -1466
rect -1596 -2410 -1572 -1490
rect -652 -2410 -628 -1490
rect -1596 -2434 -628 -2410
rect -308 -1511 12 -1469
rect -308 -2389 -266 -1511
rect -30 -2389 12 -1511
rect -308 -2431 12 -2389
rect 126 -1490 1094 -1466
rect 126 -2410 150 -1490
rect 1070 -2410 1094 -1490
rect 126 -2434 1094 -2410
rect 1414 -1511 1734 -1469
rect 1414 -2389 1456 -1511
rect 1692 -2389 1734 -1511
rect 1414 -2431 1734 -2389
rect 1848 -1490 2816 -1466
rect 1848 -2410 1872 -1490
rect 2792 -2410 2816 -1490
rect 1848 -2434 2816 -2410
rect 3136 -1511 3456 -1469
rect 3136 -2389 3178 -1511
rect 3414 -2389 3456 -1511
rect 3136 -2431 3456 -2389
rect 3570 -1490 4538 -1466
rect 3570 -2410 3594 -1490
rect 4514 -2410 4538 -1490
rect 3570 -2434 4538 -2410
rect 4858 -1511 5178 -1469
rect 4858 -2389 4900 -1511
rect 5136 -2389 5178 -1511
rect 4858 -2431 5178 -2389
rect 5292 -1490 6260 -1466
rect 5292 -2410 5316 -1490
rect 6236 -2410 6260 -1490
rect 5292 -2434 6260 -2410
rect 6580 -1511 6900 -1469
rect 6580 -2389 6622 -1511
rect 6858 -2389 6900 -1511
rect 6580 -2431 6900 -2389
rect 7014 -1490 7982 -1466
rect 7014 -2410 7038 -1490
rect 7958 -2410 7982 -1490
rect 7014 -2434 7982 -2410
rect 8302 -1511 8622 -1469
rect 8302 -2389 8344 -1511
rect 8580 -2389 8622 -1511
rect 8302 -2431 8622 -2389
rect -8160 -2766 -7840 -2434
rect -6438 -2766 -6118 -2434
rect -4716 -2766 -4396 -2434
rect -2994 -2766 -2674 -2434
rect -1272 -2766 -952 -2434
rect 450 -2766 770 -2434
rect 2172 -2766 2492 -2434
rect 3894 -2766 4214 -2434
rect 5616 -2766 5936 -2434
rect 7338 -2766 7658 -2434
rect -8484 -2790 -7516 -2766
rect -8484 -3710 -8460 -2790
rect -7540 -3710 -7516 -2790
rect -8484 -3734 -7516 -3710
rect -7196 -2811 -6876 -2769
rect -7196 -3689 -7154 -2811
rect -6918 -3689 -6876 -2811
rect -7196 -3731 -6876 -3689
rect -6762 -2790 -5794 -2766
rect -6762 -3710 -6738 -2790
rect -5818 -3710 -5794 -2790
rect -6762 -3734 -5794 -3710
rect -5474 -2811 -5154 -2769
rect -5474 -3689 -5432 -2811
rect -5196 -3689 -5154 -2811
rect -5474 -3731 -5154 -3689
rect -5040 -2790 -4072 -2766
rect -5040 -3710 -5016 -2790
rect -4096 -3710 -4072 -2790
rect -5040 -3734 -4072 -3710
rect -3752 -2811 -3432 -2769
rect -3752 -3689 -3710 -2811
rect -3474 -3689 -3432 -2811
rect -3752 -3731 -3432 -3689
rect -3318 -2790 -2350 -2766
rect -3318 -3710 -3294 -2790
rect -2374 -3710 -2350 -2790
rect -3318 -3734 -2350 -3710
rect -2030 -2811 -1710 -2769
rect -2030 -3689 -1988 -2811
rect -1752 -3689 -1710 -2811
rect -2030 -3731 -1710 -3689
rect -1596 -2790 -628 -2766
rect -1596 -3710 -1572 -2790
rect -652 -3710 -628 -2790
rect -1596 -3734 -628 -3710
rect -308 -2811 12 -2769
rect -308 -3689 -266 -2811
rect -30 -3689 12 -2811
rect -308 -3731 12 -3689
rect 126 -2790 1094 -2766
rect 126 -3710 150 -2790
rect 1070 -3710 1094 -2790
rect 126 -3734 1094 -3710
rect 1414 -2811 1734 -2769
rect 1414 -3689 1456 -2811
rect 1692 -3689 1734 -2811
rect 1414 -3731 1734 -3689
rect 1848 -2790 2816 -2766
rect 1848 -3710 1872 -2790
rect 2792 -3710 2816 -2790
rect 1848 -3734 2816 -3710
rect 3136 -2811 3456 -2769
rect 3136 -3689 3178 -2811
rect 3414 -3689 3456 -2811
rect 3136 -3731 3456 -3689
rect 3570 -2790 4538 -2766
rect 3570 -3710 3594 -2790
rect 4514 -3710 4538 -2790
rect 3570 -3734 4538 -3710
rect 4858 -2811 5178 -2769
rect 4858 -3689 4900 -2811
rect 5136 -3689 5178 -2811
rect 4858 -3731 5178 -3689
rect 5292 -2790 6260 -2766
rect 5292 -3710 5316 -2790
rect 6236 -3710 6260 -2790
rect 5292 -3734 6260 -3710
rect 6580 -2811 6900 -2769
rect 6580 -3689 6622 -2811
rect 6858 -3689 6900 -2811
rect 6580 -3731 6900 -3689
rect 7014 -2790 7982 -2766
rect 7014 -3710 7038 -2790
rect 7958 -3710 7982 -2790
rect 7014 -3734 7982 -3710
rect 8302 -2811 8622 -2769
rect 8302 -3689 8344 -2811
rect 8580 -3689 8622 -2811
rect 8302 -3731 8622 -3689
rect -8160 -3900 -7840 -3734
rect -6438 -3900 -6118 -3734
rect -4716 -3900 -4396 -3734
rect -2994 -3900 -2674 -3734
rect -1272 -3900 -952 -3734
rect 450 -3900 770 -3734
rect 2172 -3900 2492 -3734
rect 3894 -3900 4214 -3734
rect 5616 -3900 5936 -3734
rect 7338 -3900 7658 -3734
<< properties >>
string FIXED_BBOX 6898 2650 8098 3850
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 10 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
