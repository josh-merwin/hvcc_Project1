magic
tech sky130B
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -1389 1350 -1329 2550
rect -1309 1350 -1249 2550
rect -70 1350 -10 2550
rect 10 1350 70 2550
rect 1249 1350 1309 2550
rect 1329 1350 1389 2550
rect -1389 50 -1329 1250
rect -1309 50 -1249 1250
rect -70 50 -10 1250
rect 10 50 70 1250
rect 1249 50 1309 1250
rect 1329 50 1389 1250
rect -1389 -1250 -1329 -50
rect -1309 -1250 -1249 -50
rect -70 -1250 -10 -50
rect 10 -1250 70 -50
rect 1249 -1250 1309 -50
rect 1329 -1250 1389 -50
rect -1389 -2550 -1329 -1350
rect -1309 -2550 -1249 -1350
rect -70 -2550 -10 -1350
rect 10 -2550 70 -1350
rect 1249 -2550 1309 -1350
rect 1329 -2550 1389 -1350
<< metal3 >>
rect -2628 2522 -1329 2550
rect -2628 1378 -1413 2522
rect -1349 1378 -1329 2522
rect -2628 1350 -1329 1378
rect -1309 2522 -10 2550
rect -1309 1378 -94 2522
rect -30 1378 -10 2522
rect -1309 1350 -10 1378
rect 10 2522 1309 2550
rect 10 1378 1225 2522
rect 1289 1378 1309 2522
rect 10 1350 1309 1378
rect 1329 2522 2628 2550
rect 1329 1378 2544 2522
rect 2608 1378 2628 2522
rect 1329 1350 2628 1378
rect -2628 1222 -1329 1250
rect -2628 78 -1413 1222
rect -1349 78 -1329 1222
rect -2628 50 -1329 78
rect -1309 1222 -10 1250
rect -1309 78 -94 1222
rect -30 78 -10 1222
rect -1309 50 -10 78
rect 10 1222 1309 1250
rect 10 78 1225 1222
rect 1289 78 1309 1222
rect 10 50 1309 78
rect 1329 1222 2628 1250
rect 1329 78 2544 1222
rect 2608 78 2628 1222
rect 1329 50 2628 78
rect -2628 -78 -1329 -50
rect -2628 -1222 -1413 -78
rect -1349 -1222 -1329 -78
rect -2628 -1250 -1329 -1222
rect -1309 -78 -10 -50
rect -1309 -1222 -94 -78
rect -30 -1222 -10 -78
rect -1309 -1250 -10 -1222
rect 10 -78 1309 -50
rect 10 -1222 1225 -78
rect 1289 -1222 1309 -78
rect 10 -1250 1309 -1222
rect 1329 -78 2628 -50
rect 1329 -1222 2544 -78
rect 2608 -1222 2628 -78
rect 1329 -1250 2628 -1222
rect -2628 -1378 -1329 -1350
rect -2628 -2522 -1413 -1378
rect -1349 -2522 -1329 -1378
rect -2628 -2550 -1329 -2522
rect -1309 -1378 -10 -1350
rect -1309 -2522 -94 -1378
rect -30 -2522 -10 -1378
rect -1309 -2550 -10 -2522
rect 10 -1378 1309 -1350
rect 10 -2522 1225 -1378
rect 1289 -2522 1309 -1378
rect 10 -2550 1309 -2522
rect 1329 -1378 2628 -1350
rect 1329 -2522 2544 -1378
rect 2608 -2522 2628 -1378
rect 1329 -2550 2628 -2522
<< via3 >>
rect -1413 1378 -1349 2522
rect -94 1378 -30 2522
rect 1225 1378 1289 2522
rect 2544 1378 2608 2522
rect -1413 78 -1349 1222
rect -94 78 -30 1222
rect 1225 78 1289 1222
rect 2544 78 2608 1222
rect -1413 -1222 -1349 -78
rect -94 -1222 -30 -78
rect 1225 -1222 1289 -78
rect 2544 -1222 2608 -78
rect -1413 -2522 -1349 -1378
rect -94 -2522 -30 -1378
rect 1225 -2522 1289 -1378
rect 2544 -2522 2608 -1378
<< mimcap >>
rect -2528 2410 -1528 2450
rect -2528 1490 -2488 2410
rect -1568 1490 -1528 2410
rect -2528 1450 -1528 1490
rect -1209 2410 -209 2450
rect -1209 1490 -1169 2410
rect -249 1490 -209 2410
rect -1209 1450 -209 1490
rect 110 2410 1110 2450
rect 110 1490 150 2410
rect 1070 1490 1110 2410
rect 110 1450 1110 1490
rect 1429 2410 2429 2450
rect 1429 1490 1469 2410
rect 2389 1490 2429 2410
rect 1429 1450 2429 1490
rect -2528 1110 -1528 1150
rect -2528 190 -2488 1110
rect -1568 190 -1528 1110
rect -2528 150 -1528 190
rect -1209 1110 -209 1150
rect -1209 190 -1169 1110
rect -249 190 -209 1110
rect -1209 150 -209 190
rect 110 1110 1110 1150
rect 110 190 150 1110
rect 1070 190 1110 1110
rect 110 150 1110 190
rect 1429 1110 2429 1150
rect 1429 190 1469 1110
rect 2389 190 2429 1110
rect 1429 150 2429 190
rect -2528 -190 -1528 -150
rect -2528 -1110 -2488 -190
rect -1568 -1110 -1528 -190
rect -2528 -1150 -1528 -1110
rect -1209 -190 -209 -150
rect -1209 -1110 -1169 -190
rect -249 -1110 -209 -190
rect -1209 -1150 -209 -1110
rect 110 -190 1110 -150
rect 110 -1110 150 -190
rect 1070 -1110 1110 -190
rect 110 -1150 1110 -1110
rect 1429 -190 2429 -150
rect 1429 -1110 1469 -190
rect 2389 -1110 2429 -190
rect 1429 -1150 2429 -1110
rect -2528 -1490 -1528 -1450
rect -2528 -2410 -2488 -1490
rect -1568 -2410 -1528 -1490
rect -2528 -2450 -1528 -2410
rect -1209 -1490 -209 -1450
rect -1209 -2410 -1169 -1490
rect -249 -2410 -209 -1490
rect -1209 -2450 -209 -2410
rect 110 -1490 1110 -1450
rect 110 -2410 150 -1490
rect 1070 -2410 1110 -1490
rect 110 -2450 1110 -2410
rect 1429 -1490 2429 -1450
rect 1429 -2410 1469 -1490
rect 2389 -2410 2429 -1490
rect 1429 -2450 2429 -2410
<< mimcapcontact >>
rect -2488 1490 -1568 2410
rect -1169 1490 -249 2410
rect 150 1490 1070 2410
rect 1469 1490 2389 2410
rect -2488 190 -1568 1110
rect -1169 190 -249 1110
rect 150 190 1070 1110
rect 1469 190 2389 1110
rect -2488 -1110 -1568 -190
rect -1169 -1110 -249 -190
rect 150 -1110 1070 -190
rect 1469 -1110 2389 -190
rect -2488 -2410 -1568 -1490
rect -1169 -2410 -249 -1490
rect 150 -2410 1070 -1490
rect 1469 -2410 2389 -1490
<< metal4 >>
rect -2080 2411 -1976 2600
rect -1460 2538 -1356 2600
rect -1460 2522 -1333 2538
rect -2489 2410 -1567 2411
rect -2489 1490 -2488 2410
rect -1568 1490 -1567 2410
rect -2489 1489 -1567 1490
rect -2080 1111 -1976 1489
rect -1460 1378 -1413 2522
rect -1349 1378 -1333 2522
rect -761 2411 -657 2600
rect -141 2538 -37 2600
rect -141 2522 -14 2538
rect -1170 2410 -248 2411
rect -1170 1490 -1169 2410
rect -249 1490 -248 2410
rect -1170 1489 -248 1490
rect -1460 1362 -1333 1378
rect -1460 1238 -1356 1362
rect -1460 1222 -1333 1238
rect -2489 1110 -1567 1111
rect -2489 190 -2488 1110
rect -1568 190 -1567 1110
rect -2489 189 -1567 190
rect -2080 -189 -1976 189
rect -1460 78 -1413 1222
rect -1349 78 -1333 1222
rect -761 1111 -657 1489
rect -141 1378 -94 2522
rect -30 1378 -14 2522
rect 558 2411 662 2600
rect 1178 2538 1282 2600
rect 1178 2522 1305 2538
rect 149 2410 1071 2411
rect 149 1490 150 2410
rect 1070 1490 1071 2410
rect 149 1489 1071 1490
rect -141 1362 -14 1378
rect -141 1238 -37 1362
rect -141 1222 -14 1238
rect -1170 1110 -248 1111
rect -1170 190 -1169 1110
rect -249 190 -248 1110
rect -1170 189 -248 190
rect -1460 62 -1333 78
rect -1460 -62 -1356 62
rect -1460 -78 -1333 -62
rect -2489 -190 -1567 -189
rect -2489 -1110 -2488 -190
rect -1568 -1110 -1567 -190
rect -2489 -1111 -1567 -1110
rect -2080 -1489 -1976 -1111
rect -1460 -1222 -1413 -78
rect -1349 -1222 -1333 -78
rect -761 -189 -657 189
rect -141 78 -94 1222
rect -30 78 -14 1222
rect 558 1111 662 1489
rect 1178 1378 1225 2522
rect 1289 1378 1305 2522
rect 1877 2411 1981 2600
rect 2497 2538 2601 2600
rect 2497 2522 2624 2538
rect 1468 2410 2390 2411
rect 1468 1490 1469 2410
rect 2389 1490 2390 2410
rect 1468 1489 2390 1490
rect 1178 1362 1305 1378
rect 1178 1238 1282 1362
rect 1178 1222 1305 1238
rect 149 1110 1071 1111
rect 149 190 150 1110
rect 1070 190 1071 1110
rect 149 189 1071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1170 -190 -248 -189
rect -1170 -1110 -1169 -190
rect -249 -1110 -248 -190
rect -1170 -1111 -248 -1110
rect -1460 -1238 -1333 -1222
rect -1460 -1362 -1356 -1238
rect -1460 -1378 -1333 -1362
rect -2489 -1490 -1567 -1489
rect -2489 -2410 -2488 -1490
rect -1568 -2410 -1567 -1490
rect -2489 -2411 -1567 -2410
rect -2080 -2600 -1976 -2411
rect -1460 -2522 -1413 -1378
rect -1349 -2522 -1333 -1378
rect -761 -1489 -657 -1111
rect -141 -1222 -94 -78
rect -30 -1222 -14 -78
rect 558 -189 662 189
rect 1178 78 1225 1222
rect 1289 78 1305 1222
rect 1877 1111 1981 1489
rect 2497 1378 2544 2522
rect 2608 1378 2624 2522
rect 2497 1362 2624 1378
rect 2497 1238 2601 1362
rect 2497 1222 2624 1238
rect 1468 1110 2390 1111
rect 1468 190 1469 1110
rect 2389 190 2390 1110
rect 1468 189 2390 190
rect 1178 62 1305 78
rect 1178 -62 1282 62
rect 1178 -78 1305 -62
rect 149 -190 1071 -189
rect 149 -1110 150 -190
rect 1070 -1110 1071 -190
rect 149 -1111 1071 -1110
rect -141 -1238 -14 -1222
rect -141 -1362 -37 -1238
rect -141 -1378 -14 -1362
rect -1170 -1490 -248 -1489
rect -1170 -2410 -1169 -1490
rect -249 -2410 -248 -1490
rect -1170 -2411 -248 -2410
rect -1460 -2538 -1333 -2522
rect -1460 -2600 -1356 -2538
rect -761 -2600 -657 -2411
rect -141 -2522 -94 -1378
rect -30 -2522 -14 -1378
rect 558 -1489 662 -1111
rect 1178 -1222 1225 -78
rect 1289 -1222 1305 -78
rect 1877 -189 1981 189
rect 2497 78 2544 1222
rect 2608 78 2624 1222
rect 2497 62 2624 78
rect 2497 -62 2601 62
rect 2497 -78 2624 -62
rect 1468 -190 2390 -189
rect 1468 -1110 1469 -190
rect 2389 -1110 2390 -190
rect 1468 -1111 2390 -1110
rect 1178 -1238 1305 -1222
rect 1178 -1362 1282 -1238
rect 1178 -1378 1305 -1362
rect 149 -1490 1071 -1489
rect 149 -2410 150 -1490
rect 1070 -2410 1071 -1490
rect 149 -2411 1071 -2410
rect -141 -2538 -14 -2522
rect -141 -2600 -37 -2538
rect 558 -2600 662 -2411
rect 1178 -2522 1225 -1378
rect 1289 -2522 1305 -1378
rect 1877 -1489 1981 -1111
rect 2497 -1222 2544 -78
rect 2608 -1222 2624 -78
rect 2497 -1238 2624 -1222
rect 2497 -1362 2601 -1238
rect 2497 -1378 2624 -1362
rect 1468 -1490 2390 -1489
rect 1468 -2410 1469 -1490
rect 2389 -2410 2390 -1490
rect 1468 -2411 2390 -2410
rect 1178 -2538 1305 -2522
rect 1178 -2600 1282 -2538
rect 1877 -2600 1981 -2411
rect 2497 -2522 2544 -1378
rect 2608 -2522 2624 -1378
rect 2497 -2538 2624 -2522
rect 2497 -2600 2601 -2538
<< properties >>
string FIXED_BBOX 1329 1350 2529 2550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
