magic
tech sky130B
magscale 1 2
timestamp 1652200182
<< metal3 >>
rect -650 572 731 600
rect -650 -572 647 572
rect 711 -572 731 572
rect -650 -600 731 -572
<< via3 >>
rect 647 -572 711 572
<< mimcap >>
rect -550 460 450 500
rect -550 -460 -510 460
rect 410 -460 450 460
rect -550 -500 450 -460
<< mimcapcontact >>
rect -510 -460 410 460
<< metal4 >>
rect 631 572 727 701
rect -511 460 411 461
rect -511 -460 -510 460
rect 410 -460 411 460
rect -511 -461 411 -460
rect 631 -572 647 572
rect 711 -572 727 572
rect 631 -588 727 -572
<< properties >>
string FIXED_BBOX -650 -600 550 600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
