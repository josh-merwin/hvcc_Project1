magic
tech sky130B
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -2694 2434 -2674 2600
rect -2374 2434 -2354 2600
rect -2694 1134 -2674 1466
rect -2374 1134 -2354 1466
rect -2694 -166 -2674 166
rect -2374 -166 -2354 166
rect -2694 -1466 -2674 -1134
rect -2374 -1466 -2354 -1134
rect -2694 -2600 -2674 -2434
rect -2374 -2600 -2354 -2434
rect -2350 -2600 -2054 2600
rect -2030 2550 -1710 2551
rect -2030 1350 -1652 2550
rect -972 2434 -952 2600
rect -652 2434 -632 2600
rect -1596 1466 -1390 2434
rect -2030 1349 -1710 1350
rect -2030 1250 -1710 1251
rect -2030 50 -1652 1250
rect -972 1134 -952 1466
rect -652 1134 -632 1466
rect -1596 166 -1390 1134
rect -2030 49 -1710 50
rect -2030 -50 -1710 -49
rect -2030 -1250 -1652 -50
rect -972 -166 -952 166
rect -652 -166 -632 166
rect -1596 -1134 -1390 -166
rect -2030 -1251 -1710 -1250
rect -2030 -1350 -1710 -1349
rect -2030 -2550 -1652 -1350
rect -972 -1466 -952 -1134
rect -652 -1466 -632 -1134
rect -1596 -2434 -1390 -1466
rect -2030 -2551 -1710 -2550
rect -972 -2600 -952 -2434
rect -652 -2600 -632 -2434
rect -628 -2600 -332 2600
rect -308 2550 12 2551
rect -308 1350 70 2550
rect 750 2434 770 2600
rect 1070 2434 1090 2600
rect 126 1466 332 2434
rect -308 1349 12 1350
rect -308 1250 12 1251
rect -308 50 70 1250
rect 750 1134 770 1466
rect 1070 1134 1090 1466
rect 126 166 332 1134
rect -308 49 12 50
rect -308 -50 12 -49
rect -308 -1250 70 -50
rect 750 -166 770 166
rect 1070 -166 1090 166
rect 126 -1134 332 -166
rect -308 -1251 12 -1250
rect -308 -1350 12 -1349
rect -308 -2550 70 -1350
rect 750 -1466 770 -1134
rect 1070 -1466 1090 -1134
rect 126 -2434 332 -1466
rect -308 -2551 12 -2550
rect 750 -2600 770 -2434
rect 1070 -2600 1090 -2434
rect 1094 -2600 1390 2600
rect 1414 2550 1734 2551
rect 1414 1350 1792 2550
rect 2472 2434 2492 2600
rect 2792 2434 2812 2600
rect 1848 1466 2054 2434
rect 1414 1349 1734 1350
rect 1414 1250 1734 1251
rect 1414 50 1792 1250
rect 2472 1134 2492 1466
rect 2792 1134 2812 1466
rect 1848 166 2054 1134
rect 1414 49 1734 50
rect 1414 -50 1734 -49
rect 1414 -1250 1792 -50
rect 2472 -166 2492 166
rect 2792 -166 2812 166
rect 1848 -1134 2054 -166
rect 1414 -1251 1734 -1250
rect 1414 -1350 1734 -1349
rect 1414 -2550 1792 -1350
rect 2472 -1466 2492 -1134
rect 2792 -1466 2812 -1134
rect 1848 -2434 2054 -1466
rect 1414 -2551 1734 -2550
rect 2472 -2600 2492 -2434
rect 2792 -2600 2812 -2434
rect 2816 -2600 3112 2600
rect 3136 1571 3432 2551
rect 3136 1349 3456 1571
rect 3136 1029 3456 1251
rect 3136 271 3432 1029
rect 3136 49 3456 271
rect 3136 -271 3456 -49
rect 3136 -1029 3432 -271
rect 3136 -1251 3456 -1029
rect 3136 -1571 3456 -1349
rect 3136 -2551 3432 -1571
<< metal4 >>
rect -3434 2509 -1732 2550
rect -3434 1391 -1988 2509
rect -1752 1391 -1732 2509
rect -3434 1350 -1732 1391
rect -1712 2509 -10 2550
rect -1712 1391 -266 2509
rect -30 1391 -10 2509
rect -1712 1350 -10 1391
rect 10 2509 1712 2550
rect 10 1391 1456 2509
rect 1692 1391 1712 2509
rect 10 1350 1712 1391
rect 1732 2509 3434 2550
rect 1732 1391 3178 2509
rect 3414 1391 3434 2509
rect 1732 1350 3434 1391
rect -3434 1209 -1732 1250
rect -3434 91 -1988 1209
rect -1752 91 -1732 1209
rect -3434 50 -1732 91
rect -1712 1209 -10 1250
rect -1712 91 -266 1209
rect -30 91 -10 1209
rect -1712 50 -10 91
rect 10 1209 1712 1250
rect 10 91 1456 1209
rect 1692 91 1712 1209
rect 10 50 1712 91
rect 1732 1209 3434 1250
rect 1732 91 3178 1209
rect 3414 91 3434 1209
rect 1732 50 3434 91
rect -3434 -91 -1732 -50
rect -3434 -1209 -1988 -91
rect -1752 -1209 -1732 -91
rect -3434 -1250 -1732 -1209
rect -1712 -91 -10 -50
rect -1712 -1209 -266 -91
rect -30 -1209 -10 -91
rect -1712 -1250 -10 -1209
rect 10 -91 1712 -50
rect 10 -1209 1456 -91
rect 1692 -1209 1712 -91
rect 10 -1250 1712 -1209
rect 1732 -91 3434 -50
rect 1732 -1209 3178 -91
rect 3414 -1209 3434 -91
rect 1732 -1250 3434 -1209
rect -3434 -1391 -1732 -1350
rect -3434 -2509 -1988 -1391
rect -1752 -2509 -1732 -1391
rect -3434 -2550 -1732 -2509
rect -1712 -1391 -10 -1350
rect -1712 -2509 -266 -1391
rect -30 -2509 -10 -1391
rect -1712 -2550 -10 -2509
rect 10 -1391 1712 -1350
rect 10 -2509 1456 -1391
rect 1692 -2509 1712 -1391
rect 10 -2550 1712 -2509
rect 1732 -1391 3434 -1350
rect 1732 -2509 3178 -1391
rect 3414 -2509 3434 -1391
rect 1732 -2550 3434 -2509
<< via4 >>
rect -1988 1391 -1752 2509
rect -266 1391 -30 2509
rect 1456 1391 1692 2509
rect 3178 1391 3414 2509
rect -1988 91 -1752 1209
rect -266 91 -30 1209
rect 1456 91 1692 1209
rect 3178 91 3414 1209
rect -1988 -1209 -1752 -91
rect -266 -1209 -30 -91
rect 1456 -1209 1692 -91
rect 3178 -1209 3414 -91
rect -1988 -2509 -1752 -1391
rect -266 -2509 -30 -1391
rect 1456 -2509 1692 -1391
rect 3178 -2509 3414 -1391
<< mimcap2 >>
rect -3334 2410 -2334 2450
rect -3334 1490 -3294 2410
rect -2374 1490 -2334 2410
rect -3334 1450 -2334 1490
rect -1612 2410 -612 2450
rect -1612 1490 -1572 2410
rect -652 1490 -612 2410
rect -1612 1450 -612 1490
rect 110 2410 1110 2450
rect 110 1490 150 2410
rect 1070 1490 1110 2410
rect 110 1450 1110 1490
rect 1832 2410 2832 2450
rect 1832 1490 1872 2410
rect 2792 1490 2832 2410
rect 1832 1450 2832 1490
rect -3334 1110 -2334 1150
rect -3334 190 -3294 1110
rect -2374 190 -2334 1110
rect -3334 150 -2334 190
rect -1612 1110 -612 1150
rect -1612 190 -1572 1110
rect -652 190 -612 1110
rect -1612 150 -612 190
rect 110 1110 1110 1150
rect 110 190 150 1110
rect 1070 190 1110 1110
rect 110 150 1110 190
rect 1832 1110 2832 1150
rect 1832 190 1872 1110
rect 2792 190 2832 1110
rect 1832 150 2832 190
rect -3334 -190 -2334 -150
rect -3334 -1110 -3294 -190
rect -2374 -1110 -2334 -190
rect -3334 -1150 -2334 -1110
rect -1612 -190 -612 -150
rect -1612 -1110 -1572 -190
rect -652 -1110 -612 -190
rect -1612 -1150 -612 -1110
rect 110 -190 1110 -150
rect 110 -1110 150 -190
rect 1070 -1110 1110 -190
rect 110 -1150 1110 -1110
rect 1832 -190 2832 -150
rect 1832 -1110 1872 -190
rect 2792 -1110 2832 -190
rect 1832 -1150 2832 -1110
rect -3334 -1490 -2334 -1450
rect -3334 -2410 -3294 -1490
rect -2374 -2410 -2334 -1490
rect -3334 -2450 -2334 -2410
rect -1612 -1490 -612 -1450
rect -1612 -2410 -1572 -1490
rect -652 -2410 -612 -1490
rect -1612 -2450 -612 -2410
rect 110 -1490 1110 -1450
rect 110 -2410 150 -1490
rect 1070 -2410 1110 -1490
rect 110 -2450 1110 -2410
rect 1832 -1490 2832 -1450
rect 1832 -2410 1872 -1490
rect 2792 -2410 2832 -1490
rect 1832 -2450 2832 -2410
<< mimcap2contact >>
rect -3294 1490 -2374 2410
rect -1572 1490 -652 2410
rect 150 1490 1070 2410
rect 1872 1490 2792 2410
rect -3294 190 -2374 1110
rect -1572 190 -652 1110
rect 150 190 1070 1110
rect 1872 190 2792 1110
rect -3294 -1110 -2374 -190
rect -1572 -1110 -652 -190
rect 150 -1110 1070 -190
rect 1872 -1110 2792 -190
rect -3294 -2410 -2374 -1490
rect -1572 -2410 -652 -1490
rect 150 -2410 1070 -1490
rect 1872 -2410 2792 -1490
<< metal5 >>
rect -2994 2434 -2674 2600
rect -2374 2434 -2054 2600
rect -3318 2410 -2054 2434
rect -3318 1490 -3294 2410
rect -2374 1490 -2054 2410
rect -3318 1466 -2054 1490
rect -2994 1134 -2674 1466
rect -2374 1134 -2054 1466
rect -2030 2509 -1710 2551
rect -2030 1391 -1988 2509
rect -1752 1391 -1710 2509
rect -1272 2434 -952 2600
rect -652 2434 -332 2600
rect -1596 2410 -332 2434
rect -1596 1490 -1572 2410
rect -652 1490 -332 2410
rect -1596 1466 -332 1490
rect -2030 1349 -1710 1391
rect -3318 1110 -2054 1134
rect -3318 190 -3294 1110
rect -2374 190 -2054 1110
rect -3318 166 -2054 190
rect -2994 -166 -2674 166
rect -2374 -166 -2054 166
rect -2030 1209 -1710 1251
rect -2030 91 -1988 1209
rect -1752 91 -1710 1209
rect -1272 1134 -952 1466
rect -652 1134 -332 1466
rect -308 2509 12 2551
rect -308 1391 -266 2509
rect -30 1391 12 2509
rect 450 2434 770 2600
rect 1070 2434 1390 2600
rect 126 2410 1390 2434
rect 126 1490 150 2410
rect 1070 1490 1390 2410
rect 126 1466 1390 1490
rect -308 1349 12 1391
rect -1596 1110 -332 1134
rect -1596 190 -1572 1110
rect -652 190 -332 1110
rect -1596 166 -332 190
rect -2030 49 -1710 91
rect -3318 -190 -2054 -166
rect -3318 -1110 -3294 -190
rect -2374 -1110 -2054 -190
rect -3318 -1134 -2054 -1110
rect -2994 -1466 -2674 -1134
rect -2374 -1466 -2054 -1134
rect -2030 -91 -1710 -49
rect -2030 -1209 -1988 -91
rect -1752 -1209 -1710 -91
rect -1272 -166 -952 166
rect -652 -166 -332 166
rect -308 1209 12 1251
rect -308 91 -266 1209
rect -30 91 12 1209
rect 450 1134 770 1466
rect 1070 1134 1390 1466
rect 1414 2509 1734 2551
rect 1414 1391 1456 2509
rect 1692 1391 1734 2509
rect 2172 2434 2492 2600
rect 2792 2434 3112 2600
rect 1848 2410 3112 2434
rect 1848 1490 1872 2410
rect 2792 1490 3112 2410
rect 1848 1466 3112 1490
rect 1414 1349 1734 1391
rect 126 1110 1390 1134
rect 126 190 150 1110
rect 1070 190 1390 1110
rect 126 166 1390 190
rect -308 49 12 91
rect -1596 -190 -332 -166
rect -1596 -1110 -1572 -190
rect -652 -1110 -332 -190
rect -1596 -1134 -332 -1110
rect -2030 -1251 -1710 -1209
rect -3318 -1490 -2054 -1466
rect -3318 -2410 -3294 -1490
rect -2374 -2410 -2054 -1490
rect -3318 -2434 -2054 -2410
rect -2994 -2600 -2674 -2434
rect -2374 -2600 -2054 -2434
rect -2030 -1391 -1710 -1349
rect -2030 -2509 -1988 -1391
rect -1752 -2509 -1710 -1391
rect -1272 -1466 -952 -1134
rect -652 -1466 -332 -1134
rect -308 -91 12 -49
rect -308 -1209 -266 -91
rect -30 -1209 12 -91
rect 450 -166 770 166
rect 1070 -166 1390 166
rect 1414 1209 1734 1251
rect 1414 91 1456 1209
rect 1692 91 1734 1209
rect 2172 1134 2492 1466
rect 2792 1134 3112 1466
rect 3136 2509 3456 2551
rect 3136 1391 3178 2509
rect 3414 1391 3456 2509
rect 3136 1349 3456 1391
rect 1848 1110 3112 1134
rect 1848 190 1872 1110
rect 2792 190 3112 1110
rect 1848 166 3112 190
rect 1414 49 1734 91
rect 126 -190 1390 -166
rect 126 -1110 150 -190
rect 1070 -1110 1390 -190
rect 126 -1134 1390 -1110
rect -308 -1251 12 -1209
rect -1596 -1490 -332 -1466
rect -1596 -2410 -1572 -1490
rect -652 -2410 -332 -1490
rect -1596 -2434 -332 -2410
rect -2030 -2551 -1710 -2509
rect -1272 -2600 -952 -2434
rect -652 -2600 -332 -2434
rect -308 -1391 12 -1349
rect -308 -2509 -266 -1391
rect -30 -2509 12 -1391
rect 450 -1466 770 -1134
rect 1070 -1466 1390 -1134
rect 1414 -91 1734 -49
rect 1414 -1209 1456 -91
rect 1692 -1209 1734 -91
rect 2172 -166 2492 166
rect 2792 -166 3112 166
rect 3136 1209 3456 1251
rect 3136 91 3178 1209
rect 3414 91 3456 1209
rect 3136 49 3456 91
rect 1848 -190 3112 -166
rect 1848 -1110 1872 -190
rect 2792 -1110 3112 -190
rect 1848 -1134 3112 -1110
rect 1414 -1251 1734 -1209
rect 126 -1490 1390 -1466
rect 126 -2410 150 -1490
rect 1070 -2410 1390 -1490
rect 126 -2434 1390 -2410
rect -308 -2551 12 -2509
rect 450 -2600 770 -2434
rect 1070 -2600 1390 -2434
rect 1414 -1391 1734 -1349
rect 1414 -2509 1456 -1391
rect 1692 -2509 1734 -1391
rect 2172 -1466 2492 -1134
rect 2792 -1466 3112 -1134
rect 3136 -91 3456 -49
rect 3136 -1209 3178 -91
rect 3414 -1209 3456 -91
rect 3136 -1251 3456 -1209
rect 1848 -1490 3112 -1466
rect 1848 -2410 1872 -1490
rect 2792 -2410 3112 -1490
rect 1848 -2434 3112 -2410
rect 1414 -2551 1734 -2509
rect 2172 -2600 2492 -2434
rect 2792 -2600 3112 -2434
rect 3136 -1391 3456 -1349
rect 3136 -2509 3178 -1391
rect 3414 -2509 3456 -1391
rect 3136 -2551 3456 -2509
<< properties >>
string FIXED_BBOX 1732 1350 2932 2550
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
