magic
tech sky130B
magscale 1 2
timestamp 1651947127
<< pwell >>
rect -2569 -985 2569 985
<< mvnmos >>
rect -2341 527 -2241 727
rect -2183 527 -2083 727
rect -2025 527 -1925 727
rect -1867 527 -1767 727
rect -1709 527 -1609 727
rect -1551 527 -1451 727
rect -1393 527 -1293 727
rect -1235 527 -1135 727
rect -1077 527 -977 727
rect -919 527 -819 727
rect -761 527 -661 727
rect -603 527 -503 727
rect -445 527 -345 727
rect -287 527 -187 727
rect -129 527 -29 727
rect 29 527 129 727
rect 187 527 287 727
rect 345 527 445 727
rect 503 527 603 727
rect 661 527 761 727
rect 819 527 919 727
rect 977 527 1077 727
rect 1135 527 1235 727
rect 1293 527 1393 727
rect 1451 527 1551 727
rect 1609 527 1709 727
rect 1767 527 1867 727
rect 1925 527 2025 727
rect 2083 527 2183 727
rect 2241 527 2341 727
rect -2341 109 -2241 309
rect -2183 109 -2083 309
rect -2025 109 -1925 309
rect -1867 109 -1767 309
rect -1709 109 -1609 309
rect -1551 109 -1451 309
rect -1393 109 -1293 309
rect -1235 109 -1135 309
rect -1077 109 -977 309
rect -919 109 -819 309
rect -761 109 -661 309
rect -603 109 -503 309
rect -445 109 -345 309
rect -287 109 -187 309
rect -129 109 -29 309
rect 29 109 129 309
rect 187 109 287 309
rect 345 109 445 309
rect 503 109 603 309
rect 661 109 761 309
rect 819 109 919 309
rect 977 109 1077 309
rect 1135 109 1235 309
rect 1293 109 1393 309
rect 1451 109 1551 309
rect 1609 109 1709 309
rect 1767 109 1867 309
rect 1925 109 2025 309
rect 2083 109 2183 309
rect 2241 109 2341 309
rect -2341 -309 -2241 -109
rect -2183 -309 -2083 -109
rect -2025 -309 -1925 -109
rect -1867 -309 -1767 -109
rect -1709 -309 -1609 -109
rect -1551 -309 -1451 -109
rect -1393 -309 -1293 -109
rect -1235 -309 -1135 -109
rect -1077 -309 -977 -109
rect -919 -309 -819 -109
rect -761 -309 -661 -109
rect -603 -309 -503 -109
rect -445 -309 -345 -109
rect -287 -309 -187 -109
rect -129 -309 -29 -109
rect 29 -309 129 -109
rect 187 -309 287 -109
rect 345 -309 445 -109
rect 503 -309 603 -109
rect 661 -309 761 -109
rect 819 -309 919 -109
rect 977 -309 1077 -109
rect 1135 -309 1235 -109
rect 1293 -309 1393 -109
rect 1451 -309 1551 -109
rect 1609 -309 1709 -109
rect 1767 -309 1867 -109
rect 1925 -309 2025 -109
rect 2083 -309 2183 -109
rect 2241 -309 2341 -109
rect -2341 -727 -2241 -527
rect -2183 -727 -2083 -527
rect -2025 -727 -1925 -527
rect -1867 -727 -1767 -527
rect -1709 -727 -1609 -527
rect -1551 -727 -1451 -527
rect -1393 -727 -1293 -527
rect -1235 -727 -1135 -527
rect -1077 -727 -977 -527
rect -919 -727 -819 -527
rect -761 -727 -661 -527
rect -603 -727 -503 -527
rect -445 -727 -345 -527
rect -287 -727 -187 -527
rect -129 -727 -29 -527
rect 29 -727 129 -527
rect 187 -727 287 -527
rect 345 -727 445 -527
rect 503 -727 603 -527
rect 661 -727 761 -527
rect 819 -727 919 -527
rect 977 -727 1077 -527
rect 1135 -727 1235 -527
rect 1293 -727 1393 -527
rect 1451 -727 1551 -527
rect 1609 -727 1709 -527
rect 1767 -727 1867 -527
rect 1925 -727 2025 -527
rect 2083 -727 2183 -527
rect 2241 -727 2341 -527
<< mvndiff >>
rect -2399 715 -2341 727
rect -2399 539 -2387 715
rect -2353 539 -2341 715
rect -2399 527 -2341 539
rect -2241 715 -2183 727
rect -2241 539 -2229 715
rect -2195 539 -2183 715
rect -2241 527 -2183 539
rect -2083 715 -2025 727
rect -2083 539 -2071 715
rect -2037 539 -2025 715
rect -2083 527 -2025 539
rect -1925 715 -1867 727
rect -1925 539 -1913 715
rect -1879 539 -1867 715
rect -1925 527 -1867 539
rect -1767 715 -1709 727
rect -1767 539 -1755 715
rect -1721 539 -1709 715
rect -1767 527 -1709 539
rect -1609 715 -1551 727
rect -1609 539 -1597 715
rect -1563 539 -1551 715
rect -1609 527 -1551 539
rect -1451 715 -1393 727
rect -1451 539 -1439 715
rect -1405 539 -1393 715
rect -1451 527 -1393 539
rect -1293 715 -1235 727
rect -1293 539 -1281 715
rect -1247 539 -1235 715
rect -1293 527 -1235 539
rect -1135 715 -1077 727
rect -1135 539 -1123 715
rect -1089 539 -1077 715
rect -1135 527 -1077 539
rect -977 715 -919 727
rect -977 539 -965 715
rect -931 539 -919 715
rect -977 527 -919 539
rect -819 715 -761 727
rect -819 539 -807 715
rect -773 539 -761 715
rect -819 527 -761 539
rect -661 715 -603 727
rect -661 539 -649 715
rect -615 539 -603 715
rect -661 527 -603 539
rect -503 715 -445 727
rect -503 539 -491 715
rect -457 539 -445 715
rect -503 527 -445 539
rect -345 715 -287 727
rect -345 539 -333 715
rect -299 539 -287 715
rect -345 527 -287 539
rect -187 715 -129 727
rect -187 539 -175 715
rect -141 539 -129 715
rect -187 527 -129 539
rect -29 715 29 727
rect -29 539 -17 715
rect 17 539 29 715
rect -29 527 29 539
rect 129 715 187 727
rect 129 539 141 715
rect 175 539 187 715
rect 129 527 187 539
rect 287 715 345 727
rect 287 539 299 715
rect 333 539 345 715
rect 287 527 345 539
rect 445 715 503 727
rect 445 539 457 715
rect 491 539 503 715
rect 445 527 503 539
rect 603 715 661 727
rect 603 539 615 715
rect 649 539 661 715
rect 603 527 661 539
rect 761 715 819 727
rect 761 539 773 715
rect 807 539 819 715
rect 761 527 819 539
rect 919 715 977 727
rect 919 539 931 715
rect 965 539 977 715
rect 919 527 977 539
rect 1077 715 1135 727
rect 1077 539 1089 715
rect 1123 539 1135 715
rect 1077 527 1135 539
rect 1235 715 1293 727
rect 1235 539 1247 715
rect 1281 539 1293 715
rect 1235 527 1293 539
rect 1393 715 1451 727
rect 1393 539 1405 715
rect 1439 539 1451 715
rect 1393 527 1451 539
rect 1551 715 1609 727
rect 1551 539 1563 715
rect 1597 539 1609 715
rect 1551 527 1609 539
rect 1709 715 1767 727
rect 1709 539 1721 715
rect 1755 539 1767 715
rect 1709 527 1767 539
rect 1867 715 1925 727
rect 1867 539 1879 715
rect 1913 539 1925 715
rect 1867 527 1925 539
rect 2025 715 2083 727
rect 2025 539 2037 715
rect 2071 539 2083 715
rect 2025 527 2083 539
rect 2183 715 2241 727
rect 2183 539 2195 715
rect 2229 539 2241 715
rect 2183 527 2241 539
rect 2341 715 2399 727
rect 2341 539 2353 715
rect 2387 539 2399 715
rect 2341 527 2399 539
rect -2399 297 -2341 309
rect -2399 121 -2387 297
rect -2353 121 -2341 297
rect -2399 109 -2341 121
rect -2241 297 -2183 309
rect -2241 121 -2229 297
rect -2195 121 -2183 297
rect -2241 109 -2183 121
rect -2083 297 -2025 309
rect -2083 121 -2071 297
rect -2037 121 -2025 297
rect -2083 109 -2025 121
rect -1925 297 -1867 309
rect -1925 121 -1913 297
rect -1879 121 -1867 297
rect -1925 109 -1867 121
rect -1767 297 -1709 309
rect -1767 121 -1755 297
rect -1721 121 -1709 297
rect -1767 109 -1709 121
rect -1609 297 -1551 309
rect -1609 121 -1597 297
rect -1563 121 -1551 297
rect -1609 109 -1551 121
rect -1451 297 -1393 309
rect -1451 121 -1439 297
rect -1405 121 -1393 297
rect -1451 109 -1393 121
rect -1293 297 -1235 309
rect -1293 121 -1281 297
rect -1247 121 -1235 297
rect -1293 109 -1235 121
rect -1135 297 -1077 309
rect -1135 121 -1123 297
rect -1089 121 -1077 297
rect -1135 109 -1077 121
rect -977 297 -919 309
rect -977 121 -965 297
rect -931 121 -919 297
rect -977 109 -919 121
rect -819 297 -761 309
rect -819 121 -807 297
rect -773 121 -761 297
rect -819 109 -761 121
rect -661 297 -603 309
rect -661 121 -649 297
rect -615 121 -603 297
rect -661 109 -603 121
rect -503 297 -445 309
rect -503 121 -491 297
rect -457 121 -445 297
rect -503 109 -445 121
rect -345 297 -287 309
rect -345 121 -333 297
rect -299 121 -287 297
rect -345 109 -287 121
rect -187 297 -129 309
rect -187 121 -175 297
rect -141 121 -129 297
rect -187 109 -129 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 129 297 187 309
rect 129 121 141 297
rect 175 121 187 297
rect 129 109 187 121
rect 287 297 345 309
rect 287 121 299 297
rect 333 121 345 297
rect 287 109 345 121
rect 445 297 503 309
rect 445 121 457 297
rect 491 121 503 297
rect 445 109 503 121
rect 603 297 661 309
rect 603 121 615 297
rect 649 121 661 297
rect 603 109 661 121
rect 761 297 819 309
rect 761 121 773 297
rect 807 121 819 297
rect 761 109 819 121
rect 919 297 977 309
rect 919 121 931 297
rect 965 121 977 297
rect 919 109 977 121
rect 1077 297 1135 309
rect 1077 121 1089 297
rect 1123 121 1135 297
rect 1077 109 1135 121
rect 1235 297 1293 309
rect 1235 121 1247 297
rect 1281 121 1293 297
rect 1235 109 1293 121
rect 1393 297 1451 309
rect 1393 121 1405 297
rect 1439 121 1451 297
rect 1393 109 1451 121
rect 1551 297 1609 309
rect 1551 121 1563 297
rect 1597 121 1609 297
rect 1551 109 1609 121
rect 1709 297 1767 309
rect 1709 121 1721 297
rect 1755 121 1767 297
rect 1709 109 1767 121
rect 1867 297 1925 309
rect 1867 121 1879 297
rect 1913 121 1925 297
rect 1867 109 1925 121
rect 2025 297 2083 309
rect 2025 121 2037 297
rect 2071 121 2083 297
rect 2025 109 2083 121
rect 2183 297 2241 309
rect 2183 121 2195 297
rect 2229 121 2241 297
rect 2183 109 2241 121
rect 2341 297 2399 309
rect 2341 121 2353 297
rect 2387 121 2399 297
rect 2341 109 2399 121
rect -2399 -121 -2341 -109
rect -2399 -297 -2387 -121
rect -2353 -297 -2341 -121
rect -2399 -309 -2341 -297
rect -2241 -121 -2183 -109
rect -2241 -297 -2229 -121
rect -2195 -297 -2183 -121
rect -2241 -309 -2183 -297
rect -2083 -121 -2025 -109
rect -2083 -297 -2071 -121
rect -2037 -297 -2025 -121
rect -2083 -309 -2025 -297
rect -1925 -121 -1867 -109
rect -1925 -297 -1913 -121
rect -1879 -297 -1867 -121
rect -1925 -309 -1867 -297
rect -1767 -121 -1709 -109
rect -1767 -297 -1755 -121
rect -1721 -297 -1709 -121
rect -1767 -309 -1709 -297
rect -1609 -121 -1551 -109
rect -1609 -297 -1597 -121
rect -1563 -297 -1551 -121
rect -1609 -309 -1551 -297
rect -1451 -121 -1393 -109
rect -1451 -297 -1439 -121
rect -1405 -297 -1393 -121
rect -1451 -309 -1393 -297
rect -1293 -121 -1235 -109
rect -1293 -297 -1281 -121
rect -1247 -297 -1235 -121
rect -1293 -309 -1235 -297
rect -1135 -121 -1077 -109
rect -1135 -297 -1123 -121
rect -1089 -297 -1077 -121
rect -1135 -309 -1077 -297
rect -977 -121 -919 -109
rect -977 -297 -965 -121
rect -931 -297 -919 -121
rect -977 -309 -919 -297
rect -819 -121 -761 -109
rect -819 -297 -807 -121
rect -773 -297 -761 -121
rect -819 -309 -761 -297
rect -661 -121 -603 -109
rect -661 -297 -649 -121
rect -615 -297 -603 -121
rect -661 -309 -603 -297
rect -503 -121 -445 -109
rect -503 -297 -491 -121
rect -457 -297 -445 -121
rect -503 -309 -445 -297
rect -345 -121 -287 -109
rect -345 -297 -333 -121
rect -299 -297 -287 -121
rect -345 -309 -287 -297
rect -187 -121 -129 -109
rect -187 -297 -175 -121
rect -141 -297 -129 -121
rect -187 -309 -129 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 129 -121 187 -109
rect 129 -297 141 -121
rect 175 -297 187 -121
rect 129 -309 187 -297
rect 287 -121 345 -109
rect 287 -297 299 -121
rect 333 -297 345 -121
rect 287 -309 345 -297
rect 445 -121 503 -109
rect 445 -297 457 -121
rect 491 -297 503 -121
rect 445 -309 503 -297
rect 603 -121 661 -109
rect 603 -297 615 -121
rect 649 -297 661 -121
rect 603 -309 661 -297
rect 761 -121 819 -109
rect 761 -297 773 -121
rect 807 -297 819 -121
rect 761 -309 819 -297
rect 919 -121 977 -109
rect 919 -297 931 -121
rect 965 -297 977 -121
rect 919 -309 977 -297
rect 1077 -121 1135 -109
rect 1077 -297 1089 -121
rect 1123 -297 1135 -121
rect 1077 -309 1135 -297
rect 1235 -121 1293 -109
rect 1235 -297 1247 -121
rect 1281 -297 1293 -121
rect 1235 -309 1293 -297
rect 1393 -121 1451 -109
rect 1393 -297 1405 -121
rect 1439 -297 1451 -121
rect 1393 -309 1451 -297
rect 1551 -121 1609 -109
rect 1551 -297 1563 -121
rect 1597 -297 1609 -121
rect 1551 -309 1609 -297
rect 1709 -121 1767 -109
rect 1709 -297 1721 -121
rect 1755 -297 1767 -121
rect 1709 -309 1767 -297
rect 1867 -121 1925 -109
rect 1867 -297 1879 -121
rect 1913 -297 1925 -121
rect 1867 -309 1925 -297
rect 2025 -121 2083 -109
rect 2025 -297 2037 -121
rect 2071 -297 2083 -121
rect 2025 -309 2083 -297
rect 2183 -121 2241 -109
rect 2183 -297 2195 -121
rect 2229 -297 2241 -121
rect 2183 -309 2241 -297
rect 2341 -121 2399 -109
rect 2341 -297 2353 -121
rect 2387 -297 2399 -121
rect 2341 -309 2399 -297
rect -2399 -539 -2341 -527
rect -2399 -715 -2387 -539
rect -2353 -715 -2341 -539
rect -2399 -727 -2341 -715
rect -2241 -539 -2183 -527
rect -2241 -715 -2229 -539
rect -2195 -715 -2183 -539
rect -2241 -727 -2183 -715
rect -2083 -539 -2025 -527
rect -2083 -715 -2071 -539
rect -2037 -715 -2025 -539
rect -2083 -727 -2025 -715
rect -1925 -539 -1867 -527
rect -1925 -715 -1913 -539
rect -1879 -715 -1867 -539
rect -1925 -727 -1867 -715
rect -1767 -539 -1709 -527
rect -1767 -715 -1755 -539
rect -1721 -715 -1709 -539
rect -1767 -727 -1709 -715
rect -1609 -539 -1551 -527
rect -1609 -715 -1597 -539
rect -1563 -715 -1551 -539
rect -1609 -727 -1551 -715
rect -1451 -539 -1393 -527
rect -1451 -715 -1439 -539
rect -1405 -715 -1393 -539
rect -1451 -727 -1393 -715
rect -1293 -539 -1235 -527
rect -1293 -715 -1281 -539
rect -1247 -715 -1235 -539
rect -1293 -727 -1235 -715
rect -1135 -539 -1077 -527
rect -1135 -715 -1123 -539
rect -1089 -715 -1077 -539
rect -1135 -727 -1077 -715
rect -977 -539 -919 -527
rect -977 -715 -965 -539
rect -931 -715 -919 -539
rect -977 -727 -919 -715
rect -819 -539 -761 -527
rect -819 -715 -807 -539
rect -773 -715 -761 -539
rect -819 -727 -761 -715
rect -661 -539 -603 -527
rect -661 -715 -649 -539
rect -615 -715 -603 -539
rect -661 -727 -603 -715
rect -503 -539 -445 -527
rect -503 -715 -491 -539
rect -457 -715 -445 -539
rect -503 -727 -445 -715
rect -345 -539 -287 -527
rect -345 -715 -333 -539
rect -299 -715 -287 -539
rect -345 -727 -287 -715
rect -187 -539 -129 -527
rect -187 -715 -175 -539
rect -141 -715 -129 -539
rect -187 -727 -129 -715
rect -29 -539 29 -527
rect -29 -715 -17 -539
rect 17 -715 29 -539
rect -29 -727 29 -715
rect 129 -539 187 -527
rect 129 -715 141 -539
rect 175 -715 187 -539
rect 129 -727 187 -715
rect 287 -539 345 -527
rect 287 -715 299 -539
rect 333 -715 345 -539
rect 287 -727 345 -715
rect 445 -539 503 -527
rect 445 -715 457 -539
rect 491 -715 503 -539
rect 445 -727 503 -715
rect 603 -539 661 -527
rect 603 -715 615 -539
rect 649 -715 661 -539
rect 603 -727 661 -715
rect 761 -539 819 -527
rect 761 -715 773 -539
rect 807 -715 819 -539
rect 761 -727 819 -715
rect 919 -539 977 -527
rect 919 -715 931 -539
rect 965 -715 977 -539
rect 919 -727 977 -715
rect 1077 -539 1135 -527
rect 1077 -715 1089 -539
rect 1123 -715 1135 -539
rect 1077 -727 1135 -715
rect 1235 -539 1293 -527
rect 1235 -715 1247 -539
rect 1281 -715 1293 -539
rect 1235 -727 1293 -715
rect 1393 -539 1451 -527
rect 1393 -715 1405 -539
rect 1439 -715 1451 -539
rect 1393 -727 1451 -715
rect 1551 -539 1609 -527
rect 1551 -715 1563 -539
rect 1597 -715 1609 -539
rect 1551 -727 1609 -715
rect 1709 -539 1767 -527
rect 1709 -715 1721 -539
rect 1755 -715 1767 -539
rect 1709 -727 1767 -715
rect 1867 -539 1925 -527
rect 1867 -715 1879 -539
rect 1913 -715 1925 -539
rect 1867 -727 1925 -715
rect 2025 -539 2083 -527
rect 2025 -715 2037 -539
rect 2071 -715 2083 -539
rect 2025 -727 2083 -715
rect 2183 -539 2241 -527
rect 2183 -715 2195 -539
rect 2229 -715 2241 -539
rect 2183 -727 2241 -715
rect 2341 -539 2399 -527
rect 2341 -715 2353 -539
rect 2387 -715 2399 -539
rect 2341 -727 2399 -715
<< mvndiffc >>
rect -2387 539 -2353 715
rect -2229 539 -2195 715
rect -2071 539 -2037 715
rect -1913 539 -1879 715
rect -1755 539 -1721 715
rect -1597 539 -1563 715
rect -1439 539 -1405 715
rect -1281 539 -1247 715
rect -1123 539 -1089 715
rect -965 539 -931 715
rect -807 539 -773 715
rect -649 539 -615 715
rect -491 539 -457 715
rect -333 539 -299 715
rect -175 539 -141 715
rect -17 539 17 715
rect 141 539 175 715
rect 299 539 333 715
rect 457 539 491 715
rect 615 539 649 715
rect 773 539 807 715
rect 931 539 965 715
rect 1089 539 1123 715
rect 1247 539 1281 715
rect 1405 539 1439 715
rect 1563 539 1597 715
rect 1721 539 1755 715
rect 1879 539 1913 715
rect 2037 539 2071 715
rect 2195 539 2229 715
rect 2353 539 2387 715
rect -2387 121 -2353 297
rect -2229 121 -2195 297
rect -2071 121 -2037 297
rect -1913 121 -1879 297
rect -1755 121 -1721 297
rect -1597 121 -1563 297
rect -1439 121 -1405 297
rect -1281 121 -1247 297
rect -1123 121 -1089 297
rect -965 121 -931 297
rect -807 121 -773 297
rect -649 121 -615 297
rect -491 121 -457 297
rect -333 121 -299 297
rect -175 121 -141 297
rect -17 121 17 297
rect 141 121 175 297
rect 299 121 333 297
rect 457 121 491 297
rect 615 121 649 297
rect 773 121 807 297
rect 931 121 965 297
rect 1089 121 1123 297
rect 1247 121 1281 297
rect 1405 121 1439 297
rect 1563 121 1597 297
rect 1721 121 1755 297
rect 1879 121 1913 297
rect 2037 121 2071 297
rect 2195 121 2229 297
rect 2353 121 2387 297
rect -2387 -297 -2353 -121
rect -2229 -297 -2195 -121
rect -2071 -297 -2037 -121
rect -1913 -297 -1879 -121
rect -1755 -297 -1721 -121
rect -1597 -297 -1563 -121
rect -1439 -297 -1405 -121
rect -1281 -297 -1247 -121
rect -1123 -297 -1089 -121
rect -965 -297 -931 -121
rect -807 -297 -773 -121
rect -649 -297 -615 -121
rect -491 -297 -457 -121
rect -333 -297 -299 -121
rect -175 -297 -141 -121
rect -17 -297 17 -121
rect 141 -297 175 -121
rect 299 -297 333 -121
rect 457 -297 491 -121
rect 615 -297 649 -121
rect 773 -297 807 -121
rect 931 -297 965 -121
rect 1089 -297 1123 -121
rect 1247 -297 1281 -121
rect 1405 -297 1439 -121
rect 1563 -297 1597 -121
rect 1721 -297 1755 -121
rect 1879 -297 1913 -121
rect 2037 -297 2071 -121
rect 2195 -297 2229 -121
rect 2353 -297 2387 -121
rect -2387 -715 -2353 -539
rect -2229 -715 -2195 -539
rect -2071 -715 -2037 -539
rect -1913 -715 -1879 -539
rect -1755 -715 -1721 -539
rect -1597 -715 -1563 -539
rect -1439 -715 -1405 -539
rect -1281 -715 -1247 -539
rect -1123 -715 -1089 -539
rect -965 -715 -931 -539
rect -807 -715 -773 -539
rect -649 -715 -615 -539
rect -491 -715 -457 -539
rect -333 -715 -299 -539
rect -175 -715 -141 -539
rect -17 -715 17 -539
rect 141 -715 175 -539
rect 299 -715 333 -539
rect 457 -715 491 -539
rect 615 -715 649 -539
rect 773 -715 807 -539
rect 931 -715 965 -539
rect 1089 -715 1123 -539
rect 1247 -715 1281 -539
rect 1405 -715 1439 -539
rect 1563 -715 1597 -539
rect 1721 -715 1755 -539
rect 1879 -715 1913 -539
rect 2037 -715 2071 -539
rect 2195 -715 2229 -539
rect 2353 -715 2387 -539
<< mvpsubdiff >>
rect -2533 937 2533 949
rect -2533 903 -2425 937
rect 2425 903 2533 937
rect -2533 891 2533 903
rect -2533 841 -2475 891
rect -2533 -841 -2521 841
rect -2487 -841 -2475 841
rect 2475 841 2533 891
rect -2533 -891 -2475 -841
rect 2475 -841 2487 841
rect 2521 -841 2533 841
rect 2475 -891 2533 -841
rect -2533 -903 2533 -891
rect -2533 -937 -2425 -903
rect 2425 -937 2533 -903
rect -2533 -949 2533 -937
<< mvpsubdiffcont >>
rect -2425 903 2425 937
rect -2521 -841 -2487 841
rect 2487 -841 2521 841
rect -2425 -937 2425 -903
<< poly >>
rect -2341 799 -2241 815
rect -2341 765 -2325 799
rect -2257 765 -2241 799
rect -2341 727 -2241 765
rect -2183 799 -2083 815
rect -2183 765 -2167 799
rect -2099 765 -2083 799
rect -2183 727 -2083 765
rect -2025 799 -1925 815
rect -2025 765 -2009 799
rect -1941 765 -1925 799
rect -2025 727 -1925 765
rect -1867 799 -1767 815
rect -1867 765 -1851 799
rect -1783 765 -1767 799
rect -1867 727 -1767 765
rect -1709 799 -1609 815
rect -1709 765 -1693 799
rect -1625 765 -1609 799
rect -1709 727 -1609 765
rect -1551 799 -1451 815
rect -1551 765 -1535 799
rect -1467 765 -1451 799
rect -1551 727 -1451 765
rect -1393 799 -1293 815
rect -1393 765 -1377 799
rect -1309 765 -1293 799
rect -1393 727 -1293 765
rect -1235 799 -1135 815
rect -1235 765 -1219 799
rect -1151 765 -1135 799
rect -1235 727 -1135 765
rect -1077 799 -977 815
rect -1077 765 -1061 799
rect -993 765 -977 799
rect -1077 727 -977 765
rect -919 799 -819 815
rect -919 765 -903 799
rect -835 765 -819 799
rect -919 727 -819 765
rect -761 799 -661 815
rect -761 765 -745 799
rect -677 765 -661 799
rect -761 727 -661 765
rect -603 799 -503 815
rect -603 765 -587 799
rect -519 765 -503 799
rect -603 727 -503 765
rect -445 799 -345 815
rect -445 765 -429 799
rect -361 765 -345 799
rect -445 727 -345 765
rect -287 799 -187 815
rect -287 765 -271 799
rect -203 765 -187 799
rect -287 727 -187 765
rect -129 799 -29 815
rect -129 765 -113 799
rect -45 765 -29 799
rect -129 727 -29 765
rect 29 799 129 815
rect 29 765 45 799
rect 113 765 129 799
rect 29 727 129 765
rect 187 799 287 815
rect 187 765 203 799
rect 271 765 287 799
rect 187 727 287 765
rect 345 799 445 815
rect 345 765 361 799
rect 429 765 445 799
rect 345 727 445 765
rect 503 799 603 815
rect 503 765 519 799
rect 587 765 603 799
rect 503 727 603 765
rect 661 799 761 815
rect 661 765 677 799
rect 745 765 761 799
rect 661 727 761 765
rect 819 799 919 815
rect 819 765 835 799
rect 903 765 919 799
rect 819 727 919 765
rect 977 799 1077 815
rect 977 765 993 799
rect 1061 765 1077 799
rect 977 727 1077 765
rect 1135 799 1235 815
rect 1135 765 1151 799
rect 1219 765 1235 799
rect 1135 727 1235 765
rect 1293 799 1393 815
rect 1293 765 1309 799
rect 1377 765 1393 799
rect 1293 727 1393 765
rect 1451 799 1551 815
rect 1451 765 1467 799
rect 1535 765 1551 799
rect 1451 727 1551 765
rect 1609 799 1709 815
rect 1609 765 1625 799
rect 1693 765 1709 799
rect 1609 727 1709 765
rect 1767 799 1867 815
rect 1767 765 1783 799
rect 1851 765 1867 799
rect 1767 727 1867 765
rect 1925 799 2025 815
rect 1925 765 1941 799
rect 2009 765 2025 799
rect 1925 727 2025 765
rect 2083 799 2183 815
rect 2083 765 2099 799
rect 2167 765 2183 799
rect 2083 727 2183 765
rect 2241 799 2341 815
rect 2241 765 2257 799
rect 2325 765 2341 799
rect 2241 727 2341 765
rect -2341 489 -2241 527
rect -2341 455 -2325 489
rect -2257 455 -2241 489
rect -2341 439 -2241 455
rect -2183 489 -2083 527
rect -2183 455 -2167 489
rect -2099 455 -2083 489
rect -2183 439 -2083 455
rect -2025 489 -1925 527
rect -2025 455 -2009 489
rect -1941 455 -1925 489
rect -2025 439 -1925 455
rect -1867 489 -1767 527
rect -1867 455 -1851 489
rect -1783 455 -1767 489
rect -1867 439 -1767 455
rect -1709 489 -1609 527
rect -1709 455 -1693 489
rect -1625 455 -1609 489
rect -1709 439 -1609 455
rect -1551 489 -1451 527
rect -1551 455 -1535 489
rect -1467 455 -1451 489
rect -1551 439 -1451 455
rect -1393 489 -1293 527
rect -1393 455 -1377 489
rect -1309 455 -1293 489
rect -1393 439 -1293 455
rect -1235 489 -1135 527
rect -1235 455 -1219 489
rect -1151 455 -1135 489
rect -1235 439 -1135 455
rect -1077 489 -977 527
rect -1077 455 -1061 489
rect -993 455 -977 489
rect -1077 439 -977 455
rect -919 489 -819 527
rect -919 455 -903 489
rect -835 455 -819 489
rect -919 439 -819 455
rect -761 489 -661 527
rect -761 455 -745 489
rect -677 455 -661 489
rect -761 439 -661 455
rect -603 489 -503 527
rect -603 455 -587 489
rect -519 455 -503 489
rect -603 439 -503 455
rect -445 489 -345 527
rect -445 455 -429 489
rect -361 455 -345 489
rect -445 439 -345 455
rect -287 489 -187 527
rect -287 455 -271 489
rect -203 455 -187 489
rect -287 439 -187 455
rect -129 489 -29 527
rect -129 455 -113 489
rect -45 455 -29 489
rect -129 439 -29 455
rect 29 489 129 527
rect 29 455 45 489
rect 113 455 129 489
rect 29 439 129 455
rect 187 489 287 527
rect 187 455 203 489
rect 271 455 287 489
rect 187 439 287 455
rect 345 489 445 527
rect 345 455 361 489
rect 429 455 445 489
rect 345 439 445 455
rect 503 489 603 527
rect 503 455 519 489
rect 587 455 603 489
rect 503 439 603 455
rect 661 489 761 527
rect 661 455 677 489
rect 745 455 761 489
rect 661 439 761 455
rect 819 489 919 527
rect 819 455 835 489
rect 903 455 919 489
rect 819 439 919 455
rect 977 489 1077 527
rect 977 455 993 489
rect 1061 455 1077 489
rect 977 439 1077 455
rect 1135 489 1235 527
rect 1135 455 1151 489
rect 1219 455 1235 489
rect 1135 439 1235 455
rect 1293 489 1393 527
rect 1293 455 1309 489
rect 1377 455 1393 489
rect 1293 439 1393 455
rect 1451 489 1551 527
rect 1451 455 1467 489
rect 1535 455 1551 489
rect 1451 439 1551 455
rect 1609 489 1709 527
rect 1609 455 1625 489
rect 1693 455 1709 489
rect 1609 439 1709 455
rect 1767 489 1867 527
rect 1767 455 1783 489
rect 1851 455 1867 489
rect 1767 439 1867 455
rect 1925 489 2025 527
rect 1925 455 1941 489
rect 2009 455 2025 489
rect 1925 439 2025 455
rect 2083 489 2183 527
rect 2083 455 2099 489
rect 2167 455 2183 489
rect 2083 439 2183 455
rect 2241 489 2341 527
rect 2241 455 2257 489
rect 2325 455 2341 489
rect 2241 439 2341 455
rect -2341 381 -2241 397
rect -2341 347 -2325 381
rect -2257 347 -2241 381
rect -2341 309 -2241 347
rect -2183 381 -2083 397
rect -2183 347 -2167 381
rect -2099 347 -2083 381
rect -2183 309 -2083 347
rect -2025 381 -1925 397
rect -2025 347 -2009 381
rect -1941 347 -1925 381
rect -2025 309 -1925 347
rect -1867 381 -1767 397
rect -1867 347 -1851 381
rect -1783 347 -1767 381
rect -1867 309 -1767 347
rect -1709 381 -1609 397
rect -1709 347 -1693 381
rect -1625 347 -1609 381
rect -1709 309 -1609 347
rect -1551 381 -1451 397
rect -1551 347 -1535 381
rect -1467 347 -1451 381
rect -1551 309 -1451 347
rect -1393 381 -1293 397
rect -1393 347 -1377 381
rect -1309 347 -1293 381
rect -1393 309 -1293 347
rect -1235 381 -1135 397
rect -1235 347 -1219 381
rect -1151 347 -1135 381
rect -1235 309 -1135 347
rect -1077 381 -977 397
rect -1077 347 -1061 381
rect -993 347 -977 381
rect -1077 309 -977 347
rect -919 381 -819 397
rect -919 347 -903 381
rect -835 347 -819 381
rect -919 309 -819 347
rect -761 381 -661 397
rect -761 347 -745 381
rect -677 347 -661 381
rect -761 309 -661 347
rect -603 381 -503 397
rect -603 347 -587 381
rect -519 347 -503 381
rect -603 309 -503 347
rect -445 381 -345 397
rect -445 347 -429 381
rect -361 347 -345 381
rect -445 309 -345 347
rect -287 381 -187 397
rect -287 347 -271 381
rect -203 347 -187 381
rect -287 309 -187 347
rect -129 381 -29 397
rect -129 347 -113 381
rect -45 347 -29 381
rect -129 309 -29 347
rect 29 381 129 397
rect 29 347 45 381
rect 113 347 129 381
rect 29 309 129 347
rect 187 381 287 397
rect 187 347 203 381
rect 271 347 287 381
rect 187 309 287 347
rect 345 381 445 397
rect 345 347 361 381
rect 429 347 445 381
rect 345 309 445 347
rect 503 381 603 397
rect 503 347 519 381
rect 587 347 603 381
rect 503 309 603 347
rect 661 381 761 397
rect 661 347 677 381
rect 745 347 761 381
rect 661 309 761 347
rect 819 381 919 397
rect 819 347 835 381
rect 903 347 919 381
rect 819 309 919 347
rect 977 381 1077 397
rect 977 347 993 381
rect 1061 347 1077 381
rect 977 309 1077 347
rect 1135 381 1235 397
rect 1135 347 1151 381
rect 1219 347 1235 381
rect 1135 309 1235 347
rect 1293 381 1393 397
rect 1293 347 1309 381
rect 1377 347 1393 381
rect 1293 309 1393 347
rect 1451 381 1551 397
rect 1451 347 1467 381
rect 1535 347 1551 381
rect 1451 309 1551 347
rect 1609 381 1709 397
rect 1609 347 1625 381
rect 1693 347 1709 381
rect 1609 309 1709 347
rect 1767 381 1867 397
rect 1767 347 1783 381
rect 1851 347 1867 381
rect 1767 309 1867 347
rect 1925 381 2025 397
rect 1925 347 1941 381
rect 2009 347 2025 381
rect 1925 309 2025 347
rect 2083 381 2183 397
rect 2083 347 2099 381
rect 2167 347 2183 381
rect 2083 309 2183 347
rect 2241 381 2341 397
rect 2241 347 2257 381
rect 2325 347 2341 381
rect 2241 309 2341 347
rect -2341 71 -2241 109
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2341 21 -2241 37
rect -2183 71 -2083 109
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2183 21 -2083 37
rect -2025 71 -1925 109
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -2025 21 -1925 37
rect -1867 71 -1767 109
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1867 21 -1767 37
rect -1709 71 -1609 109
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1709 21 -1609 37
rect -1551 71 -1451 109
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 109
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 109
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 109
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 109
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 109
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 109
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 109
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect 1609 71 1709 109
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1609 21 1709 37
rect 1767 71 1867 109
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1767 21 1867 37
rect 1925 71 2025 109
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 1925 21 2025 37
rect 2083 71 2183 109
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2083 21 2183 37
rect 2241 71 2341 109
rect 2241 37 2257 71
rect 2325 37 2341 71
rect 2241 21 2341 37
rect -2341 -37 -2241 -21
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2341 -109 -2241 -71
rect -2183 -37 -2083 -21
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2183 -109 -2083 -71
rect -2025 -37 -1925 -21
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -2025 -109 -1925 -71
rect -1867 -37 -1767 -21
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1867 -109 -1767 -71
rect -1709 -37 -1609 -21
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1709 -109 -1609 -71
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -109 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -109 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -109 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -109 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -109 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -109 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -109 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -109 1551 -71
rect 1609 -37 1709 -21
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1609 -109 1709 -71
rect 1767 -37 1867 -21
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1767 -109 1867 -71
rect 1925 -37 2025 -21
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 1925 -109 2025 -71
rect 2083 -37 2183 -21
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2083 -109 2183 -71
rect 2241 -37 2341 -21
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect 2241 -109 2341 -71
rect -2341 -347 -2241 -309
rect -2341 -381 -2325 -347
rect -2257 -381 -2241 -347
rect -2341 -397 -2241 -381
rect -2183 -347 -2083 -309
rect -2183 -381 -2167 -347
rect -2099 -381 -2083 -347
rect -2183 -397 -2083 -381
rect -2025 -347 -1925 -309
rect -2025 -381 -2009 -347
rect -1941 -381 -1925 -347
rect -2025 -397 -1925 -381
rect -1867 -347 -1767 -309
rect -1867 -381 -1851 -347
rect -1783 -381 -1767 -347
rect -1867 -397 -1767 -381
rect -1709 -347 -1609 -309
rect -1709 -381 -1693 -347
rect -1625 -381 -1609 -347
rect -1709 -397 -1609 -381
rect -1551 -347 -1451 -309
rect -1551 -381 -1535 -347
rect -1467 -381 -1451 -347
rect -1551 -397 -1451 -381
rect -1393 -347 -1293 -309
rect -1393 -381 -1377 -347
rect -1309 -381 -1293 -347
rect -1393 -397 -1293 -381
rect -1235 -347 -1135 -309
rect -1235 -381 -1219 -347
rect -1151 -381 -1135 -347
rect -1235 -397 -1135 -381
rect -1077 -347 -977 -309
rect -1077 -381 -1061 -347
rect -993 -381 -977 -347
rect -1077 -397 -977 -381
rect -919 -347 -819 -309
rect -919 -381 -903 -347
rect -835 -381 -819 -347
rect -919 -397 -819 -381
rect -761 -347 -661 -309
rect -761 -381 -745 -347
rect -677 -381 -661 -347
rect -761 -397 -661 -381
rect -603 -347 -503 -309
rect -603 -381 -587 -347
rect -519 -381 -503 -347
rect -603 -397 -503 -381
rect -445 -347 -345 -309
rect -445 -381 -429 -347
rect -361 -381 -345 -347
rect -445 -397 -345 -381
rect -287 -347 -187 -309
rect -287 -381 -271 -347
rect -203 -381 -187 -347
rect -287 -397 -187 -381
rect -129 -347 -29 -309
rect -129 -381 -113 -347
rect -45 -381 -29 -347
rect -129 -397 -29 -381
rect 29 -347 129 -309
rect 29 -381 45 -347
rect 113 -381 129 -347
rect 29 -397 129 -381
rect 187 -347 287 -309
rect 187 -381 203 -347
rect 271 -381 287 -347
rect 187 -397 287 -381
rect 345 -347 445 -309
rect 345 -381 361 -347
rect 429 -381 445 -347
rect 345 -397 445 -381
rect 503 -347 603 -309
rect 503 -381 519 -347
rect 587 -381 603 -347
rect 503 -397 603 -381
rect 661 -347 761 -309
rect 661 -381 677 -347
rect 745 -381 761 -347
rect 661 -397 761 -381
rect 819 -347 919 -309
rect 819 -381 835 -347
rect 903 -381 919 -347
rect 819 -397 919 -381
rect 977 -347 1077 -309
rect 977 -381 993 -347
rect 1061 -381 1077 -347
rect 977 -397 1077 -381
rect 1135 -347 1235 -309
rect 1135 -381 1151 -347
rect 1219 -381 1235 -347
rect 1135 -397 1235 -381
rect 1293 -347 1393 -309
rect 1293 -381 1309 -347
rect 1377 -381 1393 -347
rect 1293 -397 1393 -381
rect 1451 -347 1551 -309
rect 1451 -381 1467 -347
rect 1535 -381 1551 -347
rect 1451 -397 1551 -381
rect 1609 -347 1709 -309
rect 1609 -381 1625 -347
rect 1693 -381 1709 -347
rect 1609 -397 1709 -381
rect 1767 -347 1867 -309
rect 1767 -381 1783 -347
rect 1851 -381 1867 -347
rect 1767 -397 1867 -381
rect 1925 -347 2025 -309
rect 1925 -381 1941 -347
rect 2009 -381 2025 -347
rect 1925 -397 2025 -381
rect 2083 -347 2183 -309
rect 2083 -381 2099 -347
rect 2167 -381 2183 -347
rect 2083 -397 2183 -381
rect 2241 -347 2341 -309
rect 2241 -381 2257 -347
rect 2325 -381 2341 -347
rect 2241 -397 2341 -381
rect -2341 -455 -2241 -439
rect -2341 -489 -2325 -455
rect -2257 -489 -2241 -455
rect -2341 -527 -2241 -489
rect -2183 -455 -2083 -439
rect -2183 -489 -2167 -455
rect -2099 -489 -2083 -455
rect -2183 -527 -2083 -489
rect -2025 -455 -1925 -439
rect -2025 -489 -2009 -455
rect -1941 -489 -1925 -455
rect -2025 -527 -1925 -489
rect -1867 -455 -1767 -439
rect -1867 -489 -1851 -455
rect -1783 -489 -1767 -455
rect -1867 -527 -1767 -489
rect -1709 -455 -1609 -439
rect -1709 -489 -1693 -455
rect -1625 -489 -1609 -455
rect -1709 -527 -1609 -489
rect -1551 -455 -1451 -439
rect -1551 -489 -1535 -455
rect -1467 -489 -1451 -455
rect -1551 -527 -1451 -489
rect -1393 -455 -1293 -439
rect -1393 -489 -1377 -455
rect -1309 -489 -1293 -455
rect -1393 -527 -1293 -489
rect -1235 -455 -1135 -439
rect -1235 -489 -1219 -455
rect -1151 -489 -1135 -455
rect -1235 -527 -1135 -489
rect -1077 -455 -977 -439
rect -1077 -489 -1061 -455
rect -993 -489 -977 -455
rect -1077 -527 -977 -489
rect -919 -455 -819 -439
rect -919 -489 -903 -455
rect -835 -489 -819 -455
rect -919 -527 -819 -489
rect -761 -455 -661 -439
rect -761 -489 -745 -455
rect -677 -489 -661 -455
rect -761 -527 -661 -489
rect -603 -455 -503 -439
rect -603 -489 -587 -455
rect -519 -489 -503 -455
rect -603 -527 -503 -489
rect -445 -455 -345 -439
rect -445 -489 -429 -455
rect -361 -489 -345 -455
rect -445 -527 -345 -489
rect -287 -455 -187 -439
rect -287 -489 -271 -455
rect -203 -489 -187 -455
rect -287 -527 -187 -489
rect -129 -455 -29 -439
rect -129 -489 -113 -455
rect -45 -489 -29 -455
rect -129 -527 -29 -489
rect 29 -455 129 -439
rect 29 -489 45 -455
rect 113 -489 129 -455
rect 29 -527 129 -489
rect 187 -455 287 -439
rect 187 -489 203 -455
rect 271 -489 287 -455
rect 187 -527 287 -489
rect 345 -455 445 -439
rect 345 -489 361 -455
rect 429 -489 445 -455
rect 345 -527 445 -489
rect 503 -455 603 -439
rect 503 -489 519 -455
rect 587 -489 603 -455
rect 503 -527 603 -489
rect 661 -455 761 -439
rect 661 -489 677 -455
rect 745 -489 761 -455
rect 661 -527 761 -489
rect 819 -455 919 -439
rect 819 -489 835 -455
rect 903 -489 919 -455
rect 819 -527 919 -489
rect 977 -455 1077 -439
rect 977 -489 993 -455
rect 1061 -489 1077 -455
rect 977 -527 1077 -489
rect 1135 -455 1235 -439
rect 1135 -489 1151 -455
rect 1219 -489 1235 -455
rect 1135 -527 1235 -489
rect 1293 -455 1393 -439
rect 1293 -489 1309 -455
rect 1377 -489 1393 -455
rect 1293 -527 1393 -489
rect 1451 -455 1551 -439
rect 1451 -489 1467 -455
rect 1535 -489 1551 -455
rect 1451 -527 1551 -489
rect 1609 -455 1709 -439
rect 1609 -489 1625 -455
rect 1693 -489 1709 -455
rect 1609 -527 1709 -489
rect 1767 -455 1867 -439
rect 1767 -489 1783 -455
rect 1851 -489 1867 -455
rect 1767 -527 1867 -489
rect 1925 -455 2025 -439
rect 1925 -489 1941 -455
rect 2009 -489 2025 -455
rect 1925 -527 2025 -489
rect 2083 -455 2183 -439
rect 2083 -489 2099 -455
rect 2167 -489 2183 -455
rect 2083 -527 2183 -489
rect 2241 -455 2341 -439
rect 2241 -489 2257 -455
rect 2325 -489 2341 -455
rect 2241 -527 2341 -489
rect -2341 -765 -2241 -727
rect -2341 -799 -2325 -765
rect -2257 -799 -2241 -765
rect -2341 -815 -2241 -799
rect -2183 -765 -2083 -727
rect -2183 -799 -2167 -765
rect -2099 -799 -2083 -765
rect -2183 -815 -2083 -799
rect -2025 -765 -1925 -727
rect -2025 -799 -2009 -765
rect -1941 -799 -1925 -765
rect -2025 -815 -1925 -799
rect -1867 -765 -1767 -727
rect -1867 -799 -1851 -765
rect -1783 -799 -1767 -765
rect -1867 -815 -1767 -799
rect -1709 -765 -1609 -727
rect -1709 -799 -1693 -765
rect -1625 -799 -1609 -765
rect -1709 -815 -1609 -799
rect -1551 -765 -1451 -727
rect -1551 -799 -1535 -765
rect -1467 -799 -1451 -765
rect -1551 -815 -1451 -799
rect -1393 -765 -1293 -727
rect -1393 -799 -1377 -765
rect -1309 -799 -1293 -765
rect -1393 -815 -1293 -799
rect -1235 -765 -1135 -727
rect -1235 -799 -1219 -765
rect -1151 -799 -1135 -765
rect -1235 -815 -1135 -799
rect -1077 -765 -977 -727
rect -1077 -799 -1061 -765
rect -993 -799 -977 -765
rect -1077 -815 -977 -799
rect -919 -765 -819 -727
rect -919 -799 -903 -765
rect -835 -799 -819 -765
rect -919 -815 -819 -799
rect -761 -765 -661 -727
rect -761 -799 -745 -765
rect -677 -799 -661 -765
rect -761 -815 -661 -799
rect -603 -765 -503 -727
rect -603 -799 -587 -765
rect -519 -799 -503 -765
rect -603 -815 -503 -799
rect -445 -765 -345 -727
rect -445 -799 -429 -765
rect -361 -799 -345 -765
rect -445 -815 -345 -799
rect -287 -765 -187 -727
rect -287 -799 -271 -765
rect -203 -799 -187 -765
rect -287 -815 -187 -799
rect -129 -765 -29 -727
rect -129 -799 -113 -765
rect -45 -799 -29 -765
rect -129 -815 -29 -799
rect 29 -765 129 -727
rect 29 -799 45 -765
rect 113 -799 129 -765
rect 29 -815 129 -799
rect 187 -765 287 -727
rect 187 -799 203 -765
rect 271 -799 287 -765
rect 187 -815 287 -799
rect 345 -765 445 -727
rect 345 -799 361 -765
rect 429 -799 445 -765
rect 345 -815 445 -799
rect 503 -765 603 -727
rect 503 -799 519 -765
rect 587 -799 603 -765
rect 503 -815 603 -799
rect 661 -765 761 -727
rect 661 -799 677 -765
rect 745 -799 761 -765
rect 661 -815 761 -799
rect 819 -765 919 -727
rect 819 -799 835 -765
rect 903 -799 919 -765
rect 819 -815 919 -799
rect 977 -765 1077 -727
rect 977 -799 993 -765
rect 1061 -799 1077 -765
rect 977 -815 1077 -799
rect 1135 -765 1235 -727
rect 1135 -799 1151 -765
rect 1219 -799 1235 -765
rect 1135 -815 1235 -799
rect 1293 -765 1393 -727
rect 1293 -799 1309 -765
rect 1377 -799 1393 -765
rect 1293 -815 1393 -799
rect 1451 -765 1551 -727
rect 1451 -799 1467 -765
rect 1535 -799 1551 -765
rect 1451 -815 1551 -799
rect 1609 -765 1709 -727
rect 1609 -799 1625 -765
rect 1693 -799 1709 -765
rect 1609 -815 1709 -799
rect 1767 -765 1867 -727
rect 1767 -799 1783 -765
rect 1851 -799 1867 -765
rect 1767 -815 1867 -799
rect 1925 -765 2025 -727
rect 1925 -799 1941 -765
rect 2009 -799 2025 -765
rect 1925 -815 2025 -799
rect 2083 -765 2183 -727
rect 2083 -799 2099 -765
rect 2167 -799 2183 -765
rect 2083 -815 2183 -799
rect 2241 -765 2341 -727
rect 2241 -799 2257 -765
rect 2325 -799 2341 -765
rect 2241 -815 2341 -799
<< polycont >>
rect -2325 765 -2257 799
rect -2167 765 -2099 799
rect -2009 765 -1941 799
rect -1851 765 -1783 799
rect -1693 765 -1625 799
rect -1535 765 -1467 799
rect -1377 765 -1309 799
rect -1219 765 -1151 799
rect -1061 765 -993 799
rect -903 765 -835 799
rect -745 765 -677 799
rect -587 765 -519 799
rect -429 765 -361 799
rect -271 765 -203 799
rect -113 765 -45 799
rect 45 765 113 799
rect 203 765 271 799
rect 361 765 429 799
rect 519 765 587 799
rect 677 765 745 799
rect 835 765 903 799
rect 993 765 1061 799
rect 1151 765 1219 799
rect 1309 765 1377 799
rect 1467 765 1535 799
rect 1625 765 1693 799
rect 1783 765 1851 799
rect 1941 765 2009 799
rect 2099 765 2167 799
rect 2257 765 2325 799
rect -2325 455 -2257 489
rect -2167 455 -2099 489
rect -2009 455 -1941 489
rect -1851 455 -1783 489
rect -1693 455 -1625 489
rect -1535 455 -1467 489
rect -1377 455 -1309 489
rect -1219 455 -1151 489
rect -1061 455 -993 489
rect -903 455 -835 489
rect -745 455 -677 489
rect -587 455 -519 489
rect -429 455 -361 489
rect -271 455 -203 489
rect -113 455 -45 489
rect 45 455 113 489
rect 203 455 271 489
rect 361 455 429 489
rect 519 455 587 489
rect 677 455 745 489
rect 835 455 903 489
rect 993 455 1061 489
rect 1151 455 1219 489
rect 1309 455 1377 489
rect 1467 455 1535 489
rect 1625 455 1693 489
rect 1783 455 1851 489
rect 1941 455 2009 489
rect 2099 455 2167 489
rect 2257 455 2325 489
rect -2325 347 -2257 381
rect -2167 347 -2099 381
rect -2009 347 -1941 381
rect -1851 347 -1783 381
rect -1693 347 -1625 381
rect -1535 347 -1467 381
rect -1377 347 -1309 381
rect -1219 347 -1151 381
rect -1061 347 -993 381
rect -903 347 -835 381
rect -745 347 -677 381
rect -587 347 -519 381
rect -429 347 -361 381
rect -271 347 -203 381
rect -113 347 -45 381
rect 45 347 113 381
rect 203 347 271 381
rect 361 347 429 381
rect 519 347 587 381
rect 677 347 745 381
rect 835 347 903 381
rect 993 347 1061 381
rect 1151 347 1219 381
rect 1309 347 1377 381
rect 1467 347 1535 381
rect 1625 347 1693 381
rect 1783 347 1851 381
rect 1941 347 2009 381
rect 2099 347 2167 381
rect 2257 347 2325 381
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect -2325 -381 -2257 -347
rect -2167 -381 -2099 -347
rect -2009 -381 -1941 -347
rect -1851 -381 -1783 -347
rect -1693 -381 -1625 -347
rect -1535 -381 -1467 -347
rect -1377 -381 -1309 -347
rect -1219 -381 -1151 -347
rect -1061 -381 -993 -347
rect -903 -381 -835 -347
rect -745 -381 -677 -347
rect -587 -381 -519 -347
rect -429 -381 -361 -347
rect -271 -381 -203 -347
rect -113 -381 -45 -347
rect 45 -381 113 -347
rect 203 -381 271 -347
rect 361 -381 429 -347
rect 519 -381 587 -347
rect 677 -381 745 -347
rect 835 -381 903 -347
rect 993 -381 1061 -347
rect 1151 -381 1219 -347
rect 1309 -381 1377 -347
rect 1467 -381 1535 -347
rect 1625 -381 1693 -347
rect 1783 -381 1851 -347
rect 1941 -381 2009 -347
rect 2099 -381 2167 -347
rect 2257 -381 2325 -347
rect -2325 -489 -2257 -455
rect -2167 -489 -2099 -455
rect -2009 -489 -1941 -455
rect -1851 -489 -1783 -455
rect -1693 -489 -1625 -455
rect -1535 -489 -1467 -455
rect -1377 -489 -1309 -455
rect -1219 -489 -1151 -455
rect -1061 -489 -993 -455
rect -903 -489 -835 -455
rect -745 -489 -677 -455
rect -587 -489 -519 -455
rect -429 -489 -361 -455
rect -271 -489 -203 -455
rect -113 -489 -45 -455
rect 45 -489 113 -455
rect 203 -489 271 -455
rect 361 -489 429 -455
rect 519 -489 587 -455
rect 677 -489 745 -455
rect 835 -489 903 -455
rect 993 -489 1061 -455
rect 1151 -489 1219 -455
rect 1309 -489 1377 -455
rect 1467 -489 1535 -455
rect 1625 -489 1693 -455
rect 1783 -489 1851 -455
rect 1941 -489 2009 -455
rect 2099 -489 2167 -455
rect 2257 -489 2325 -455
rect -2325 -799 -2257 -765
rect -2167 -799 -2099 -765
rect -2009 -799 -1941 -765
rect -1851 -799 -1783 -765
rect -1693 -799 -1625 -765
rect -1535 -799 -1467 -765
rect -1377 -799 -1309 -765
rect -1219 -799 -1151 -765
rect -1061 -799 -993 -765
rect -903 -799 -835 -765
rect -745 -799 -677 -765
rect -587 -799 -519 -765
rect -429 -799 -361 -765
rect -271 -799 -203 -765
rect -113 -799 -45 -765
rect 45 -799 113 -765
rect 203 -799 271 -765
rect 361 -799 429 -765
rect 519 -799 587 -765
rect 677 -799 745 -765
rect 835 -799 903 -765
rect 993 -799 1061 -765
rect 1151 -799 1219 -765
rect 1309 -799 1377 -765
rect 1467 -799 1535 -765
rect 1625 -799 1693 -765
rect 1783 -799 1851 -765
rect 1941 -799 2009 -765
rect 2099 -799 2167 -765
rect 2257 -799 2325 -765
<< locali >>
rect -2521 903 -2425 937
rect 2425 903 2521 937
rect -2521 841 -2487 903
rect 2487 841 2521 903
rect -2341 765 -2325 799
rect -2257 765 -2241 799
rect -2183 765 -2167 799
rect -2099 765 -2083 799
rect -2025 765 -2009 799
rect -1941 765 -1925 799
rect -1867 765 -1851 799
rect -1783 765 -1767 799
rect -1709 765 -1693 799
rect -1625 765 -1609 799
rect -1551 765 -1535 799
rect -1467 765 -1451 799
rect -1393 765 -1377 799
rect -1309 765 -1293 799
rect -1235 765 -1219 799
rect -1151 765 -1135 799
rect -1077 765 -1061 799
rect -993 765 -977 799
rect -919 765 -903 799
rect -835 765 -819 799
rect -761 765 -745 799
rect -677 765 -661 799
rect -603 765 -587 799
rect -519 765 -503 799
rect -445 765 -429 799
rect -361 765 -345 799
rect -287 765 -271 799
rect -203 765 -187 799
rect -129 765 -113 799
rect -45 765 -29 799
rect 29 765 45 799
rect 113 765 129 799
rect 187 765 203 799
rect 271 765 287 799
rect 345 765 361 799
rect 429 765 445 799
rect 503 765 519 799
rect 587 765 603 799
rect 661 765 677 799
rect 745 765 761 799
rect 819 765 835 799
rect 903 765 919 799
rect 977 765 993 799
rect 1061 765 1077 799
rect 1135 765 1151 799
rect 1219 765 1235 799
rect 1293 765 1309 799
rect 1377 765 1393 799
rect 1451 765 1467 799
rect 1535 765 1551 799
rect 1609 765 1625 799
rect 1693 765 1709 799
rect 1767 765 1783 799
rect 1851 765 1867 799
rect 1925 765 1941 799
rect 2009 765 2025 799
rect 2083 765 2099 799
rect 2167 765 2183 799
rect 2241 765 2257 799
rect 2325 765 2341 799
rect -2387 715 -2353 731
rect -2387 523 -2353 539
rect -2229 715 -2195 731
rect -2229 523 -2195 539
rect -2071 715 -2037 731
rect -2071 523 -2037 539
rect -1913 715 -1879 731
rect -1913 523 -1879 539
rect -1755 715 -1721 731
rect -1755 523 -1721 539
rect -1597 715 -1563 731
rect -1597 523 -1563 539
rect -1439 715 -1405 731
rect -1439 523 -1405 539
rect -1281 715 -1247 731
rect -1281 523 -1247 539
rect -1123 715 -1089 731
rect -1123 523 -1089 539
rect -965 715 -931 731
rect -965 523 -931 539
rect -807 715 -773 731
rect -807 523 -773 539
rect -649 715 -615 731
rect -649 523 -615 539
rect -491 715 -457 731
rect -491 523 -457 539
rect -333 715 -299 731
rect -333 523 -299 539
rect -175 715 -141 731
rect -175 523 -141 539
rect -17 715 17 731
rect -17 523 17 539
rect 141 715 175 731
rect 141 523 175 539
rect 299 715 333 731
rect 299 523 333 539
rect 457 715 491 731
rect 457 523 491 539
rect 615 715 649 731
rect 615 523 649 539
rect 773 715 807 731
rect 773 523 807 539
rect 931 715 965 731
rect 931 523 965 539
rect 1089 715 1123 731
rect 1089 523 1123 539
rect 1247 715 1281 731
rect 1247 523 1281 539
rect 1405 715 1439 731
rect 1405 523 1439 539
rect 1563 715 1597 731
rect 1563 523 1597 539
rect 1721 715 1755 731
rect 1721 523 1755 539
rect 1879 715 1913 731
rect 1879 523 1913 539
rect 2037 715 2071 731
rect 2037 523 2071 539
rect 2195 715 2229 731
rect 2195 523 2229 539
rect 2353 715 2387 731
rect 2353 523 2387 539
rect -2341 455 -2325 489
rect -2257 455 -2241 489
rect -2183 455 -2167 489
rect -2099 455 -2083 489
rect -2025 455 -2009 489
rect -1941 455 -1925 489
rect -1867 455 -1851 489
rect -1783 455 -1767 489
rect -1709 455 -1693 489
rect -1625 455 -1609 489
rect -1551 455 -1535 489
rect -1467 455 -1451 489
rect -1393 455 -1377 489
rect -1309 455 -1293 489
rect -1235 455 -1219 489
rect -1151 455 -1135 489
rect -1077 455 -1061 489
rect -993 455 -977 489
rect -919 455 -903 489
rect -835 455 -819 489
rect -761 455 -745 489
rect -677 455 -661 489
rect -603 455 -587 489
rect -519 455 -503 489
rect -445 455 -429 489
rect -361 455 -345 489
rect -287 455 -271 489
rect -203 455 -187 489
rect -129 455 -113 489
rect -45 455 -29 489
rect 29 455 45 489
rect 113 455 129 489
rect 187 455 203 489
rect 271 455 287 489
rect 345 455 361 489
rect 429 455 445 489
rect 503 455 519 489
rect 587 455 603 489
rect 661 455 677 489
rect 745 455 761 489
rect 819 455 835 489
rect 903 455 919 489
rect 977 455 993 489
rect 1061 455 1077 489
rect 1135 455 1151 489
rect 1219 455 1235 489
rect 1293 455 1309 489
rect 1377 455 1393 489
rect 1451 455 1467 489
rect 1535 455 1551 489
rect 1609 455 1625 489
rect 1693 455 1709 489
rect 1767 455 1783 489
rect 1851 455 1867 489
rect 1925 455 1941 489
rect 2009 455 2025 489
rect 2083 455 2099 489
rect 2167 455 2183 489
rect 2241 455 2257 489
rect 2325 455 2341 489
rect -2341 347 -2325 381
rect -2257 347 -2241 381
rect -2183 347 -2167 381
rect -2099 347 -2083 381
rect -2025 347 -2009 381
rect -1941 347 -1925 381
rect -1867 347 -1851 381
rect -1783 347 -1767 381
rect -1709 347 -1693 381
rect -1625 347 -1609 381
rect -1551 347 -1535 381
rect -1467 347 -1451 381
rect -1393 347 -1377 381
rect -1309 347 -1293 381
rect -1235 347 -1219 381
rect -1151 347 -1135 381
rect -1077 347 -1061 381
rect -993 347 -977 381
rect -919 347 -903 381
rect -835 347 -819 381
rect -761 347 -745 381
rect -677 347 -661 381
rect -603 347 -587 381
rect -519 347 -503 381
rect -445 347 -429 381
rect -361 347 -345 381
rect -287 347 -271 381
rect -203 347 -187 381
rect -129 347 -113 381
rect -45 347 -29 381
rect 29 347 45 381
rect 113 347 129 381
rect 187 347 203 381
rect 271 347 287 381
rect 345 347 361 381
rect 429 347 445 381
rect 503 347 519 381
rect 587 347 603 381
rect 661 347 677 381
rect 745 347 761 381
rect 819 347 835 381
rect 903 347 919 381
rect 977 347 993 381
rect 1061 347 1077 381
rect 1135 347 1151 381
rect 1219 347 1235 381
rect 1293 347 1309 381
rect 1377 347 1393 381
rect 1451 347 1467 381
rect 1535 347 1551 381
rect 1609 347 1625 381
rect 1693 347 1709 381
rect 1767 347 1783 381
rect 1851 347 1867 381
rect 1925 347 1941 381
rect 2009 347 2025 381
rect 2083 347 2099 381
rect 2167 347 2183 381
rect 2241 347 2257 381
rect 2325 347 2341 381
rect -2387 297 -2353 313
rect -2387 105 -2353 121
rect -2229 297 -2195 313
rect -2229 105 -2195 121
rect -2071 297 -2037 313
rect -2071 105 -2037 121
rect -1913 297 -1879 313
rect -1913 105 -1879 121
rect -1755 297 -1721 313
rect -1755 105 -1721 121
rect -1597 297 -1563 313
rect -1597 105 -1563 121
rect -1439 297 -1405 313
rect -1439 105 -1405 121
rect -1281 297 -1247 313
rect -1281 105 -1247 121
rect -1123 297 -1089 313
rect -1123 105 -1089 121
rect -965 297 -931 313
rect -965 105 -931 121
rect -807 297 -773 313
rect -807 105 -773 121
rect -649 297 -615 313
rect -649 105 -615 121
rect -491 297 -457 313
rect -491 105 -457 121
rect -333 297 -299 313
rect -333 105 -299 121
rect -175 297 -141 313
rect -175 105 -141 121
rect -17 297 17 313
rect -17 105 17 121
rect 141 297 175 313
rect 141 105 175 121
rect 299 297 333 313
rect 299 105 333 121
rect 457 297 491 313
rect 457 105 491 121
rect 615 297 649 313
rect 615 105 649 121
rect 773 297 807 313
rect 773 105 807 121
rect 931 297 965 313
rect 931 105 965 121
rect 1089 297 1123 313
rect 1089 105 1123 121
rect 1247 297 1281 313
rect 1247 105 1281 121
rect 1405 297 1439 313
rect 1405 105 1439 121
rect 1563 297 1597 313
rect 1563 105 1597 121
rect 1721 297 1755 313
rect 1721 105 1755 121
rect 1879 297 1913 313
rect 1879 105 1913 121
rect 2037 297 2071 313
rect 2037 105 2071 121
rect 2195 297 2229 313
rect 2195 105 2229 121
rect 2353 297 2387 313
rect 2353 105 2387 121
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2241 37 2257 71
rect 2325 37 2341 71
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect -2387 -121 -2353 -105
rect -2387 -313 -2353 -297
rect -2229 -121 -2195 -105
rect -2229 -313 -2195 -297
rect -2071 -121 -2037 -105
rect -2071 -313 -2037 -297
rect -1913 -121 -1879 -105
rect -1913 -313 -1879 -297
rect -1755 -121 -1721 -105
rect -1755 -313 -1721 -297
rect -1597 -121 -1563 -105
rect -1597 -313 -1563 -297
rect -1439 -121 -1405 -105
rect -1439 -313 -1405 -297
rect -1281 -121 -1247 -105
rect -1281 -313 -1247 -297
rect -1123 -121 -1089 -105
rect -1123 -313 -1089 -297
rect -965 -121 -931 -105
rect -965 -313 -931 -297
rect -807 -121 -773 -105
rect -807 -313 -773 -297
rect -649 -121 -615 -105
rect -649 -313 -615 -297
rect -491 -121 -457 -105
rect -491 -313 -457 -297
rect -333 -121 -299 -105
rect -333 -313 -299 -297
rect -175 -121 -141 -105
rect -175 -313 -141 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 141 -121 175 -105
rect 141 -313 175 -297
rect 299 -121 333 -105
rect 299 -313 333 -297
rect 457 -121 491 -105
rect 457 -313 491 -297
rect 615 -121 649 -105
rect 615 -313 649 -297
rect 773 -121 807 -105
rect 773 -313 807 -297
rect 931 -121 965 -105
rect 931 -313 965 -297
rect 1089 -121 1123 -105
rect 1089 -313 1123 -297
rect 1247 -121 1281 -105
rect 1247 -313 1281 -297
rect 1405 -121 1439 -105
rect 1405 -313 1439 -297
rect 1563 -121 1597 -105
rect 1563 -313 1597 -297
rect 1721 -121 1755 -105
rect 1721 -313 1755 -297
rect 1879 -121 1913 -105
rect 1879 -313 1913 -297
rect 2037 -121 2071 -105
rect 2037 -313 2071 -297
rect 2195 -121 2229 -105
rect 2195 -313 2229 -297
rect 2353 -121 2387 -105
rect 2353 -313 2387 -297
rect -2341 -381 -2325 -347
rect -2257 -381 -2241 -347
rect -2183 -381 -2167 -347
rect -2099 -381 -2083 -347
rect -2025 -381 -2009 -347
rect -1941 -381 -1925 -347
rect -1867 -381 -1851 -347
rect -1783 -381 -1767 -347
rect -1709 -381 -1693 -347
rect -1625 -381 -1609 -347
rect -1551 -381 -1535 -347
rect -1467 -381 -1451 -347
rect -1393 -381 -1377 -347
rect -1309 -381 -1293 -347
rect -1235 -381 -1219 -347
rect -1151 -381 -1135 -347
rect -1077 -381 -1061 -347
rect -993 -381 -977 -347
rect -919 -381 -903 -347
rect -835 -381 -819 -347
rect -761 -381 -745 -347
rect -677 -381 -661 -347
rect -603 -381 -587 -347
rect -519 -381 -503 -347
rect -445 -381 -429 -347
rect -361 -381 -345 -347
rect -287 -381 -271 -347
rect -203 -381 -187 -347
rect -129 -381 -113 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 113 -381 129 -347
rect 187 -381 203 -347
rect 271 -381 287 -347
rect 345 -381 361 -347
rect 429 -381 445 -347
rect 503 -381 519 -347
rect 587 -381 603 -347
rect 661 -381 677 -347
rect 745 -381 761 -347
rect 819 -381 835 -347
rect 903 -381 919 -347
rect 977 -381 993 -347
rect 1061 -381 1077 -347
rect 1135 -381 1151 -347
rect 1219 -381 1235 -347
rect 1293 -381 1309 -347
rect 1377 -381 1393 -347
rect 1451 -381 1467 -347
rect 1535 -381 1551 -347
rect 1609 -381 1625 -347
rect 1693 -381 1709 -347
rect 1767 -381 1783 -347
rect 1851 -381 1867 -347
rect 1925 -381 1941 -347
rect 2009 -381 2025 -347
rect 2083 -381 2099 -347
rect 2167 -381 2183 -347
rect 2241 -381 2257 -347
rect 2325 -381 2341 -347
rect -2341 -489 -2325 -455
rect -2257 -489 -2241 -455
rect -2183 -489 -2167 -455
rect -2099 -489 -2083 -455
rect -2025 -489 -2009 -455
rect -1941 -489 -1925 -455
rect -1867 -489 -1851 -455
rect -1783 -489 -1767 -455
rect -1709 -489 -1693 -455
rect -1625 -489 -1609 -455
rect -1551 -489 -1535 -455
rect -1467 -489 -1451 -455
rect -1393 -489 -1377 -455
rect -1309 -489 -1293 -455
rect -1235 -489 -1219 -455
rect -1151 -489 -1135 -455
rect -1077 -489 -1061 -455
rect -993 -489 -977 -455
rect -919 -489 -903 -455
rect -835 -489 -819 -455
rect -761 -489 -745 -455
rect -677 -489 -661 -455
rect -603 -489 -587 -455
rect -519 -489 -503 -455
rect -445 -489 -429 -455
rect -361 -489 -345 -455
rect -287 -489 -271 -455
rect -203 -489 -187 -455
rect -129 -489 -113 -455
rect -45 -489 -29 -455
rect 29 -489 45 -455
rect 113 -489 129 -455
rect 187 -489 203 -455
rect 271 -489 287 -455
rect 345 -489 361 -455
rect 429 -489 445 -455
rect 503 -489 519 -455
rect 587 -489 603 -455
rect 661 -489 677 -455
rect 745 -489 761 -455
rect 819 -489 835 -455
rect 903 -489 919 -455
rect 977 -489 993 -455
rect 1061 -489 1077 -455
rect 1135 -489 1151 -455
rect 1219 -489 1235 -455
rect 1293 -489 1309 -455
rect 1377 -489 1393 -455
rect 1451 -489 1467 -455
rect 1535 -489 1551 -455
rect 1609 -489 1625 -455
rect 1693 -489 1709 -455
rect 1767 -489 1783 -455
rect 1851 -489 1867 -455
rect 1925 -489 1941 -455
rect 2009 -489 2025 -455
rect 2083 -489 2099 -455
rect 2167 -489 2183 -455
rect 2241 -489 2257 -455
rect 2325 -489 2341 -455
rect -2387 -539 -2353 -523
rect -2387 -731 -2353 -715
rect -2229 -539 -2195 -523
rect -2229 -731 -2195 -715
rect -2071 -539 -2037 -523
rect -2071 -731 -2037 -715
rect -1913 -539 -1879 -523
rect -1913 -731 -1879 -715
rect -1755 -539 -1721 -523
rect -1755 -731 -1721 -715
rect -1597 -539 -1563 -523
rect -1597 -731 -1563 -715
rect -1439 -539 -1405 -523
rect -1439 -731 -1405 -715
rect -1281 -539 -1247 -523
rect -1281 -731 -1247 -715
rect -1123 -539 -1089 -523
rect -1123 -731 -1089 -715
rect -965 -539 -931 -523
rect -965 -731 -931 -715
rect -807 -539 -773 -523
rect -807 -731 -773 -715
rect -649 -539 -615 -523
rect -649 -731 -615 -715
rect -491 -539 -457 -523
rect -491 -731 -457 -715
rect -333 -539 -299 -523
rect -333 -731 -299 -715
rect -175 -539 -141 -523
rect -175 -731 -141 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 141 -539 175 -523
rect 141 -731 175 -715
rect 299 -539 333 -523
rect 299 -731 333 -715
rect 457 -539 491 -523
rect 457 -731 491 -715
rect 615 -539 649 -523
rect 615 -731 649 -715
rect 773 -539 807 -523
rect 773 -731 807 -715
rect 931 -539 965 -523
rect 931 -731 965 -715
rect 1089 -539 1123 -523
rect 1089 -731 1123 -715
rect 1247 -539 1281 -523
rect 1247 -731 1281 -715
rect 1405 -539 1439 -523
rect 1405 -731 1439 -715
rect 1563 -539 1597 -523
rect 1563 -731 1597 -715
rect 1721 -539 1755 -523
rect 1721 -731 1755 -715
rect 1879 -539 1913 -523
rect 1879 -731 1913 -715
rect 2037 -539 2071 -523
rect 2037 -731 2071 -715
rect 2195 -539 2229 -523
rect 2195 -731 2229 -715
rect 2353 -539 2387 -523
rect 2353 -731 2387 -715
rect -2341 -799 -2325 -765
rect -2257 -799 -2241 -765
rect -2183 -799 -2167 -765
rect -2099 -799 -2083 -765
rect -2025 -799 -2009 -765
rect -1941 -799 -1925 -765
rect -1867 -799 -1851 -765
rect -1783 -799 -1767 -765
rect -1709 -799 -1693 -765
rect -1625 -799 -1609 -765
rect -1551 -799 -1535 -765
rect -1467 -799 -1451 -765
rect -1393 -799 -1377 -765
rect -1309 -799 -1293 -765
rect -1235 -799 -1219 -765
rect -1151 -799 -1135 -765
rect -1077 -799 -1061 -765
rect -993 -799 -977 -765
rect -919 -799 -903 -765
rect -835 -799 -819 -765
rect -761 -799 -745 -765
rect -677 -799 -661 -765
rect -603 -799 -587 -765
rect -519 -799 -503 -765
rect -445 -799 -429 -765
rect -361 -799 -345 -765
rect -287 -799 -271 -765
rect -203 -799 -187 -765
rect -129 -799 -113 -765
rect -45 -799 -29 -765
rect 29 -799 45 -765
rect 113 -799 129 -765
rect 187 -799 203 -765
rect 271 -799 287 -765
rect 345 -799 361 -765
rect 429 -799 445 -765
rect 503 -799 519 -765
rect 587 -799 603 -765
rect 661 -799 677 -765
rect 745 -799 761 -765
rect 819 -799 835 -765
rect 903 -799 919 -765
rect 977 -799 993 -765
rect 1061 -799 1077 -765
rect 1135 -799 1151 -765
rect 1219 -799 1235 -765
rect 1293 -799 1309 -765
rect 1377 -799 1393 -765
rect 1451 -799 1467 -765
rect 1535 -799 1551 -765
rect 1609 -799 1625 -765
rect 1693 -799 1709 -765
rect 1767 -799 1783 -765
rect 1851 -799 1867 -765
rect 1925 -799 1941 -765
rect 2009 -799 2025 -765
rect 2083 -799 2099 -765
rect 2167 -799 2183 -765
rect 2241 -799 2257 -765
rect 2325 -799 2341 -765
rect -2521 -903 -2487 -841
rect 2487 -903 2521 -841
rect -2521 -937 -2425 -903
rect 2425 -937 2521 -903
<< viali >>
rect -2325 765 -2257 799
rect -2167 765 -2099 799
rect -2009 765 -1941 799
rect -1851 765 -1783 799
rect -1693 765 -1625 799
rect -1535 765 -1467 799
rect -1377 765 -1309 799
rect -1219 765 -1151 799
rect -1061 765 -993 799
rect -903 765 -835 799
rect -745 765 -677 799
rect -587 765 -519 799
rect -429 765 -361 799
rect -271 765 -203 799
rect -113 765 -45 799
rect 45 765 113 799
rect 203 765 271 799
rect 361 765 429 799
rect 519 765 587 799
rect 677 765 745 799
rect 835 765 903 799
rect 993 765 1061 799
rect 1151 765 1219 799
rect 1309 765 1377 799
rect 1467 765 1535 799
rect 1625 765 1693 799
rect 1783 765 1851 799
rect 1941 765 2009 799
rect 2099 765 2167 799
rect 2257 765 2325 799
rect -2387 539 -2353 715
rect -2229 539 -2195 715
rect -2071 539 -2037 715
rect -1913 539 -1879 715
rect -1755 539 -1721 715
rect -1597 539 -1563 715
rect -1439 539 -1405 715
rect -1281 539 -1247 715
rect -1123 539 -1089 715
rect -965 539 -931 715
rect -807 539 -773 715
rect -649 539 -615 715
rect -491 539 -457 715
rect -333 539 -299 715
rect -175 539 -141 715
rect -17 539 17 715
rect 141 539 175 715
rect 299 539 333 715
rect 457 539 491 715
rect 615 539 649 715
rect 773 539 807 715
rect 931 539 965 715
rect 1089 539 1123 715
rect 1247 539 1281 715
rect 1405 539 1439 715
rect 1563 539 1597 715
rect 1721 539 1755 715
rect 1879 539 1913 715
rect 2037 539 2071 715
rect 2195 539 2229 715
rect 2353 539 2387 715
rect -2325 455 -2257 489
rect -2167 455 -2099 489
rect -2009 455 -1941 489
rect -1851 455 -1783 489
rect -1693 455 -1625 489
rect -1535 455 -1467 489
rect -1377 455 -1309 489
rect -1219 455 -1151 489
rect -1061 455 -993 489
rect -903 455 -835 489
rect -745 455 -677 489
rect -587 455 -519 489
rect -429 455 -361 489
rect -271 455 -203 489
rect -113 455 -45 489
rect 45 455 113 489
rect 203 455 271 489
rect 361 455 429 489
rect 519 455 587 489
rect 677 455 745 489
rect 835 455 903 489
rect 993 455 1061 489
rect 1151 455 1219 489
rect 1309 455 1377 489
rect 1467 455 1535 489
rect 1625 455 1693 489
rect 1783 455 1851 489
rect 1941 455 2009 489
rect 2099 455 2167 489
rect 2257 455 2325 489
rect -2325 347 -2257 381
rect -2167 347 -2099 381
rect -2009 347 -1941 381
rect -1851 347 -1783 381
rect -1693 347 -1625 381
rect -1535 347 -1467 381
rect -1377 347 -1309 381
rect -1219 347 -1151 381
rect -1061 347 -993 381
rect -903 347 -835 381
rect -745 347 -677 381
rect -587 347 -519 381
rect -429 347 -361 381
rect -271 347 -203 381
rect -113 347 -45 381
rect 45 347 113 381
rect 203 347 271 381
rect 361 347 429 381
rect 519 347 587 381
rect 677 347 745 381
rect 835 347 903 381
rect 993 347 1061 381
rect 1151 347 1219 381
rect 1309 347 1377 381
rect 1467 347 1535 381
rect 1625 347 1693 381
rect 1783 347 1851 381
rect 1941 347 2009 381
rect 2099 347 2167 381
rect 2257 347 2325 381
rect -2387 121 -2353 297
rect -2229 121 -2195 297
rect -2071 121 -2037 297
rect -1913 121 -1879 297
rect -1755 121 -1721 297
rect -1597 121 -1563 297
rect -1439 121 -1405 297
rect -1281 121 -1247 297
rect -1123 121 -1089 297
rect -965 121 -931 297
rect -807 121 -773 297
rect -649 121 -615 297
rect -491 121 -457 297
rect -333 121 -299 297
rect -175 121 -141 297
rect -17 121 17 297
rect 141 121 175 297
rect 299 121 333 297
rect 457 121 491 297
rect 615 121 649 297
rect 773 121 807 297
rect 931 121 965 297
rect 1089 121 1123 297
rect 1247 121 1281 297
rect 1405 121 1439 297
rect 1563 121 1597 297
rect 1721 121 1755 297
rect 1879 121 1913 297
rect 2037 121 2071 297
rect 2195 121 2229 297
rect 2353 121 2387 297
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect -2387 -297 -2353 -121
rect -2229 -297 -2195 -121
rect -2071 -297 -2037 -121
rect -1913 -297 -1879 -121
rect -1755 -297 -1721 -121
rect -1597 -297 -1563 -121
rect -1439 -297 -1405 -121
rect -1281 -297 -1247 -121
rect -1123 -297 -1089 -121
rect -965 -297 -931 -121
rect -807 -297 -773 -121
rect -649 -297 -615 -121
rect -491 -297 -457 -121
rect -333 -297 -299 -121
rect -175 -297 -141 -121
rect -17 -297 17 -121
rect 141 -297 175 -121
rect 299 -297 333 -121
rect 457 -297 491 -121
rect 615 -297 649 -121
rect 773 -297 807 -121
rect 931 -297 965 -121
rect 1089 -297 1123 -121
rect 1247 -297 1281 -121
rect 1405 -297 1439 -121
rect 1563 -297 1597 -121
rect 1721 -297 1755 -121
rect 1879 -297 1913 -121
rect 2037 -297 2071 -121
rect 2195 -297 2229 -121
rect 2353 -297 2387 -121
rect -2325 -381 -2257 -347
rect -2167 -381 -2099 -347
rect -2009 -381 -1941 -347
rect -1851 -381 -1783 -347
rect -1693 -381 -1625 -347
rect -1535 -381 -1467 -347
rect -1377 -381 -1309 -347
rect -1219 -381 -1151 -347
rect -1061 -381 -993 -347
rect -903 -381 -835 -347
rect -745 -381 -677 -347
rect -587 -381 -519 -347
rect -429 -381 -361 -347
rect -271 -381 -203 -347
rect -113 -381 -45 -347
rect 45 -381 113 -347
rect 203 -381 271 -347
rect 361 -381 429 -347
rect 519 -381 587 -347
rect 677 -381 745 -347
rect 835 -381 903 -347
rect 993 -381 1061 -347
rect 1151 -381 1219 -347
rect 1309 -381 1377 -347
rect 1467 -381 1535 -347
rect 1625 -381 1693 -347
rect 1783 -381 1851 -347
rect 1941 -381 2009 -347
rect 2099 -381 2167 -347
rect 2257 -381 2325 -347
rect -2325 -489 -2257 -455
rect -2167 -489 -2099 -455
rect -2009 -489 -1941 -455
rect -1851 -489 -1783 -455
rect -1693 -489 -1625 -455
rect -1535 -489 -1467 -455
rect -1377 -489 -1309 -455
rect -1219 -489 -1151 -455
rect -1061 -489 -993 -455
rect -903 -489 -835 -455
rect -745 -489 -677 -455
rect -587 -489 -519 -455
rect -429 -489 -361 -455
rect -271 -489 -203 -455
rect -113 -489 -45 -455
rect 45 -489 113 -455
rect 203 -489 271 -455
rect 361 -489 429 -455
rect 519 -489 587 -455
rect 677 -489 745 -455
rect 835 -489 903 -455
rect 993 -489 1061 -455
rect 1151 -489 1219 -455
rect 1309 -489 1377 -455
rect 1467 -489 1535 -455
rect 1625 -489 1693 -455
rect 1783 -489 1851 -455
rect 1941 -489 2009 -455
rect 2099 -489 2167 -455
rect 2257 -489 2325 -455
rect -2387 -715 -2353 -539
rect -2229 -715 -2195 -539
rect -2071 -715 -2037 -539
rect -1913 -715 -1879 -539
rect -1755 -715 -1721 -539
rect -1597 -715 -1563 -539
rect -1439 -715 -1405 -539
rect -1281 -715 -1247 -539
rect -1123 -715 -1089 -539
rect -965 -715 -931 -539
rect -807 -715 -773 -539
rect -649 -715 -615 -539
rect -491 -715 -457 -539
rect -333 -715 -299 -539
rect -175 -715 -141 -539
rect -17 -715 17 -539
rect 141 -715 175 -539
rect 299 -715 333 -539
rect 457 -715 491 -539
rect 615 -715 649 -539
rect 773 -715 807 -539
rect 931 -715 965 -539
rect 1089 -715 1123 -539
rect 1247 -715 1281 -539
rect 1405 -715 1439 -539
rect 1563 -715 1597 -539
rect 1721 -715 1755 -539
rect 1879 -715 1913 -539
rect 2037 -715 2071 -539
rect 2195 -715 2229 -539
rect 2353 -715 2387 -539
rect -2325 -799 -2257 -765
rect -2167 -799 -2099 -765
rect -2009 -799 -1941 -765
rect -1851 -799 -1783 -765
rect -1693 -799 -1625 -765
rect -1535 -799 -1467 -765
rect -1377 -799 -1309 -765
rect -1219 -799 -1151 -765
rect -1061 -799 -993 -765
rect -903 -799 -835 -765
rect -745 -799 -677 -765
rect -587 -799 -519 -765
rect -429 -799 -361 -765
rect -271 -799 -203 -765
rect -113 -799 -45 -765
rect 45 -799 113 -765
rect 203 -799 271 -765
rect 361 -799 429 -765
rect 519 -799 587 -765
rect 677 -799 745 -765
rect 835 -799 903 -765
rect 993 -799 1061 -765
rect 1151 -799 1219 -765
rect 1309 -799 1377 -765
rect 1467 -799 1535 -765
rect 1625 -799 1693 -765
rect 1783 -799 1851 -765
rect 1941 -799 2009 -765
rect 2099 -799 2167 -765
rect 2257 -799 2325 -765
<< metal1 >>
rect -2337 799 -2245 805
rect -2337 765 -2325 799
rect -2257 765 -2245 799
rect -2337 759 -2245 765
rect -2179 799 -2087 805
rect -2179 765 -2167 799
rect -2099 765 -2087 799
rect -2179 759 -2087 765
rect -2021 799 -1929 805
rect -2021 765 -2009 799
rect -1941 765 -1929 799
rect -2021 759 -1929 765
rect -1863 799 -1771 805
rect -1863 765 -1851 799
rect -1783 765 -1771 799
rect -1863 759 -1771 765
rect -1705 799 -1613 805
rect -1705 765 -1693 799
rect -1625 765 -1613 799
rect -1705 759 -1613 765
rect -1547 799 -1455 805
rect -1547 765 -1535 799
rect -1467 765 -1455 799
rect -1547 759 -1455 765
rect -1389 799 -1297 805
rect -1389 765 -1377 799
rect -1309 765 -1297 799
rect -1389 759 -1297 765
rect -1231 799 -1139 805
rect -1231 765 -1219 799
rect -1151 765 -1139 799
rect -1231 759 -1139 765
rect -1073 799 -981 805
rect -1073 765 -1061 799
rect -993 765 -981 799
rect -1073 759 -981 765
rect -915 799 -823 805
rect -915 765 -903 799
rect -835 765 -823 799
rect -915 759 -823 765
rect -757 799 -665 805
rect -757 765 -745 799
rect -677 765 -665 799
rect -757 759 -665 765
rect -599 799 -507 805
rect -599 765 -587 799
rect -519 765 -507 799
rect -599 759 -507 765
rect -441 799 -349 805
rect -441 765 -429 799
rect -361 765 -349 799
rect -441 759 -349 765
rect -283 799 -191 805
rect -283 765 -271 799
rect -203 765 -191 799
rect -283 759 -191 765
rect -125 799 -33 805
rect -125 765 -113 799
rect -45 765 -33 799
rect -125 759 -33 765
rect 33 799 125 805
rect 33 765 45 799
rect 113 765 125 799
rect 33 759 125 765
rect 191 799 283 805
rect 191 765 203 799
rect 271 765 283 799
rect 191 759 283 765
rect 349 799 441 805
rect 349 765 361 799
rect 429 765 441 799
rect 349 759 441 765
rect 507 799 599 805
rect 507 765 519 799
rect 587 765 599 799
rect 507 759 599 765
rect 665 799 757 805
rect 665 765 677 799
rect 745 765 757 799
rect 665 759 757 765
rect 823 799 915 805
rect 823 765 835 799
rect 903 765 915 799
rect 823 759 915 765
rect 981 799 1073 805
rect 981 765 993 799
rect 1061 765 1073 799
rect 981 759 1073 765
rect 1139 799 1231 805
rect 1139 765 1151 799
rect 1219 765 1231 799
rect 1139 759 1231 765
rect 1297 799 1389 805
rect 1297 765 1309 799
rect 1377 765 1389 799
rect 1297 759 1389 765
rect 1455 799 1547 805
rect 1455 765 1467 799
rect 1535 765 1547 799
rect 1455 759 1547 765
rect 1613 799 1705 805
rect 1613 765 1625 799
rect 1693 765 1705 799
rect 1613 759 1705 765
rect 1771 799 1863 805
rect 1771 765 1783 799
rect 1851 765 1863 799
rect 1771 759 1863 765
rect 1929 799 2021 805
rect 1929 765 1941 799
rect 2009 765 2021 799
rect 1929 759 2021 765
rect 2087 799 2179 805
rect 2087 765 2099 799
rect 2167 765 2179 799
rect 2087 759 2179 765
rect 2245 799 2337 805
rect 2245 765 2257 799
rect 2325 765 2337 799
rect 2245 759 2337 765
rect -2393 715 -2347 727
rect -2393 539 -2387 715
rect -2353 539 -2347 715
rect -2393 527 -2347 539
rect -2235 715 -2189 727
rect -2235 539 -2229 715
rect -2195 539 -2189 715
rect -2235 527 -2189 539
rect -2077 715 -2031 727
rect -2077 539 -2071 715
rect -2037 539 -2031 715
rect -2077 527 -2031 539
rect -1919 715 -1873 727
rect -1919 539 -1913 715
rect -1879 539 -1873 715
rect -1919 527 -1873 539
rect -1761 715 -1715 727
rect -1761 539 -1755 715
rect -1721 539 -1715 715
rect -1761 527 -1715 539
rect -1603 715 -1557 727
rect -1603 539 -1597 715
rect -1563 539 -1557 715
rect -1603 527 -1557 539
rect -1445 715 -1399 727
rect -1445 539 -1439 715
rect -1405 539 -1399 715
rect -1445 527 -1399 539
rect -1287 715 -1241 727
rect -1287 539 -1281 715
rect -1247 539 -1241 715
rect -1287 527 -1241 539
rect -1129 715 -1083 727
rect -1129 539 -1123 715
rect -1089 539 -1083 715
rect -1129 527 -1083 539
rect -971 715 -925 727
rect -971 539 -965 715
rect -931 539 -925 715
rect -971 527 -925 539
rect -813 715 -767 727
rect -813 539 -807 715
rect -773 539 -767 715
rect -813 527 -767 539
rect -655 715 -609 727
rect -655 539 -649 715
rect -615 539 -609 715
rect -655 527 -609 539
rect -497 715 -451 727
rect -497 539 -491 715
rect -457 539 -451 715
rect -497 527 -451 539
rect -339 715 -293 727
rect -339 539 -333 715
rect -299 539 -293 715
rect -339 527 -293 539
rect -181 715 -135 727
rect -181 539 -175 715
rect -141 539 -135 715
rect -181 527 -135 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 135 715 181 727
rect 135 539 141 715
rect 175 539 181 715
rect 135 527 181 539
rect 293 715 339 727
rect 293 539 299 715
rect 333 539 339 715
rect 293 527 339 539
rect 451 715 497 727
rect 451 539 457 715
rect 491 539 497 715
rect 451 527 497 539
rect 609 715 655 727
rect 609 539 615 715
rect 649 539 655 715
rect 609 527 655 539
rect 767 715 813 727
rect 767 539 773 715
rect 807 539 813 715
rect 767 527 813 539
rect 925 715 971 727
rect 925 539 931 715
rect 965 539 971 715
rect 925 527 971 539
rect 1083 715 1129 727
rect 1083 539 1089 715
rect 1123 539 1129 715
rect 1083 527 1129 539
rect 1241 715 1287 727
rect 1241 539 1247 715
rect 1281 539 1287 715
rect 1241 527 1287 539
rect 1399 715 1445 727
rect 1399 539 1405 715
rect 1439 539 1445 715
rect 1399 527 1445 539
rect 1557 715 1603 727
rect 1557 539 1563 715
rect 1597 539 1603 715
rect 1557 527 1603 539
rect 1715 715 1761 727
rect 1715 539 1721 715
rect 1755 539 1761 715
rect 1715 527 1761 539
rect 1873 715 1919 727
rect 1873 539 1879 715
rect 1913 539 1919 715
rect 1873 527 1919 539
rect 2031 715 2077 727
rect 2031 539 2037 715
rect 2071 539 2077 715
rect 2031 527 2077 539
rect 2189 715 2235 727
rect 2189 539 2195 715
rect 2229 539 2235 715
rect 2189 527 2235 539
rect 2347 715 2393 727
rect 2347 539 2353 715
rect 2387 539 2393 715
rect 2347 527 2393 539
rect -2337 489 -2245 495
rect -2337 455 -2325 489
rect -2257 455 -2245 489
rect -2337 449 -2245 455
rect -2179 489 -2087 495
rect -2179 455 -2167 489
rect -2099 455 -2087 489
rect -2179 449 -2087 455
rect -2021 489 -1929 495
rect -2021 455 -2009 489
rect -1941 455 -1929 489
rect -2021 449 -1929 455
rect -1863 489 -1771 495
rect -1863 455 -1851 489
rect -1783 455 -1771 489
rect -1863 449 -1771 455
rect -1705 489 -1613 495
rect -1705 455 -1693 489
rect -1625 455 -1613 489
rect -1705 449 -1613 455
rect -1547 489 -1455 495
rect -1547 455 -1535 489
rect -1467 455 -1455 489
rect -1547 449 -1455 455
rect -1389 489 -1297 495
rect -1389 455 -1377 489
rect -1309 455 -1297 489
rect -1389 449 -1297 455
rect -1231 489 -1139 495
rect -1231 455 -1219 489
rect -1151 455 -1139 489
rect -1231 449 -1139 455
rect -1073 489 -981 495
rect -1073 455 -1061 489
rect -993 455 -981 489
rect -1073 449 -981 455
rect -915 489 -823 495
rect -915 455 -903 489
rect -835 455 -823 489
rect -915 449 -823 455
rect -757 489 -665 495
rect -757 455 -745 489
rect -677 455 -665 489
rect -757 449 -665 455
rect -599 489 -507 495
rect -599 455 -587 489
rect -519 455 -507 489
rect -599 449 -507 455
rect -441 489 -349 495
rect -441 455 -429 489
rect -361 455 -349 489
rect -441 449 -349 455
rect -283 489 -191 495
rect -283 455 -271 489
rect -203 455 -191 489
rect -283 449 -191 455
rect -125 489 -33 495
rect -125 455 -113 489
rect -45 455 -33 489
rect -125 449 -33 455
rect 33 489 125 495
rect 33 455 45 489
rect 113 455 125 489
rect 33 449 125 455
rect 191 489 283 495
rect 191 455 203 489
rect 271 455 283 489
rect 191 449 283 455
rect 349 489 441 495
rect 349 455 361 489
rect 429 455 441 489
rect 349 449 441 455
rect 507 489 599 495
rect 507 455 519 489
rect 587 455 599 489
rect 507 449 599 455
rect 665 489 757 495
rect 665 455 677 489
rect 745 455 757 489
rect 665 449 757 455
rect 823 489 915 495
rect 823 455 835 489
rect 903 455 915 489
rect 823 449 915 455
rect 981 489 1073 495
rect 981 455 993 489
rect 1061 455 1073 489
rect 981 449 1073 455
rect 1139 489 1231 495
rect 1139 455 1151 489
rect 1219 455 1231 489
rect 1139 449 1231 455
rect 1297 489 1389 495
rect 1297 455 1309 489
rect 1377 455 1389 489
rect 1297 449 1389 455
rect 1455 489 1547 495
rect 1455 455 1467 489
rect 1535 455 1547 489
rect 1455 449 1547 455
rect 1613 489 1705 495
rect 1613 455 1625 489
rect 1693 455 1705 489
rect 1613 449 1705 455
rect 1771 489 1863 495
rect 1771 455 1783 489
rect 1851 455 1863 489
rect 1771 449 1863 455
rect 1929 489 2021 495
rect 1929 455 1941 489
rect 2009 455 2021 489
rect 1929 449 2021 455
rect 2087 489 2179 495
rect 2087 455 2099 489
rect 2167 455 2179 489
rect 2087 449 2179 455
rect 2245 489 2337 495
rect 2245 455 2257 489
rect 2325 455 2337 489
rect 2245 449 2337 455
rect -2337 381 -2245 387
rect -2337 347 -2325 381
rect -2257 347 -2245 381
rect -2337 341 -2245 347
rect -2179 381 -2087 387
rect -2179 347 -2167 381
rect -2099 347 -2087 381
rect -2179 341 -2087 347
rect -2021 381 -1929 387
rect -2021 347 -2009 381
rect -1941 347 -1929 381
rect -2021 341 -1929 347
rect -1863 381 -1771 387
rect -1863 347 -1851 381
rect -1783 347 -1771 381
rect -1863 341 -1771 347
rect -1705 381 -1613 387
rect -1705 347 -1693 381
rect -1625 347 -1613 381
rect -1705 341 -1613 347
rect -1547 381 -1455 387
rect -1547 347 -1535 381
rect -1467 347 -1455 381
rect -1547 341 -1455 347
rect -1389 381 -1297 387
rect -1389 347 -1377 381
rect -1309 347 -1297 381
rect -1389 341 -1297 347
rect -1231 381 -1139 387
rect -1231 347 -1219 381
rect -1151 347 -1139 381
rect -1231 341 -1139 347
rect -1073 381 -981 387
rect -1073 347 -1061 381
rect -993 347 -981 381
rect -1073 341 -981 347
rect -915 381 -823 387
rect -915 347 -903 381
rect -835 347 -823 381
rect -915 341 -823 347
rect -757 381 -665 387
rect -757 347 -745 381
rect -677 347 -665 381
rect -757 341 -665 347
rect -599 381 -507 387
rect -599 347 -587 381
rect -519 347 -507 381
rect -599 341 -507 347
rect -441 381 -349 387
rect -441 347 -429 381
rect -361 347 -349 381
rect -441 341 -349 347
rect -283 381 -191 387
rect -283 347 -271 381
rect -203 347 -191 381
rect -283 341 -191 347
rect -125 381 -33 387
rect -125 347 -113 381
rect -45 347 -33 381
rect -125 341 -33 347
rect 33 381 125 387
rect 33 347 45 381
rect 113 347 125 381
rect 33 341 125 347
rect 191 381 283 387
rect 191 347 203 381
rect 271 347 283 381
rect 191 341 283 347
rect 349 381 441 387
rect 349 347 361 381
rect 429 347 441 381
rect 349 341 441 347
rect 507 381 599 387
rect 507 347 519 381
rect 587 347 599 381
rect 507 341 599 347
rect 665 381 757 387
rect 665 347 677 381
rect 745 347 757 381
rect 665 341 757 347
rect 823 381 915 387
rect 823 347 835 381
rect 903 347 915 381
rect 823 341 915 347
rect 981 381 1073 387
rect 981 347 993 381
rect 1061 347 1073 381
rect 981 341 1073 347
rect 1139 381 1231 387
rect 1139 347 1151 381
rect 1219 347 1231 381
rect 1139 341 1231 347
rect 1297 381 1389 387
rect 1297 347 1309 381
rect 1377 347 1389 381
rect 1297 341 1389 347
rect 1455 381 1547 387
rect 1455 347 1467 381
rect 1535 347 1547 381
rect 1455 341 1547 347
rect 1613 381 1705 387
rect 1613 347 1625 381
rect 1693 347 1705 381
rect 1613 341 1705 347
rect 1771 381 1863 387
rect 1771 347 1783 381
rect 1851 347 1863 381
rect 1771 341 1863 347
rect 1929 381 2021 387
rect 1929 347 1941 381
rect 2009 347 2021 381
rect 1929 341 2021 347
rect 2087 381 2179 387
rect 2087 347 2099 381
rect 2167 347 2179 381
rect 2087 341 2179 347
rect 2245 381 2337 387
rect 2245 347 2257 381
rect 2325 347 2337 381
rect 2245 341 2337 347
rect -2393 297 -2347 309
rect -2393 121 -2387 297
rect -2353 121 -2347 297
rect -2393 109 -2347 121
rect -2235 297 -2189 309
rect -2235 121 -2229 297
rect -2195 121 -2189 297
rect -2235 109 -2189 121
rect -2077 297 -2031 309
rect -2077 121 -2071 297
rect -2037 121 -2031 297
rect -2077 109 -2031 121
rect -1919 297 -1873 309
rect -1919 121 -1913 297
rect -1879 121 -1873 297
rect -1919 109 -1873 121
rect -1761 297 -1715 309
rect -1761 121 -1755 297
rect -1721 121 -1715 297
rect -1761 109 -1715 121
rect -1603 297 -1557 309
rect -1603 121 -1597 297
rect -1563 121 -1557 297
rect -1603 109 -1557 121
rect -1445 297 -1399 309
rect -1445 121 -1439 297
rect -1405 121 -1399 297
rect -1445 109 -1399 121
rect -1287 297 -1241 309
rect -1287 121 -1281 297
rect -1247 121 -1241 297
rect -1287 109 -1241 121
rect -1129 297 -1083 309
rect -1129 121 -1123 297
rect -1089 121 -1083 297
rect -1129 109 -1083 121
rect -971 297 -925 309
rect -971 121 -965 297
rect -931 121 -925 297
rect -971 109 -925 121
rect -813 297 -767 309
rect -813 121 -807 297
rect -773 121 -767 297
rect -813 109 -767 121
rect -655 297 -609 309
rect -655 121 -649 297
rect -615 121 -609 297
rect -655 109 -609 121
rect -497 297 -451 309
rect -497 121 -491 297
rect -457 121 -451 297
rect -497 109 -451 121
rect -339 297 -293 309
rect -339 121 -333 297
rect -299 121 -293 297
rect -339 109 -293 121
rect -181 297 -135 309
rect -181 121 -175 297
rect -141 121 -135 297
rect -181 109 -135 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 135 297 181 309
rect 135 121 141 297
rect 175 121 181 297
rect 135 109 181 121
rect 293 297 339 309
rect 293 121 299 297
rect 333 121 339 297
rect 293 109 339 121
rect 451 297 497 309
rect 451 121 457 297
rect 491 121 497 297
rect 451 109 497 121
rect 609 297 655 309
rect 609 121 615 297
rect 649 121 655 297
rect 609 109 655 121
rect 767 297 813 309
rect 767 121 773 297
rect 807 121 813 297
rect 767 109 813 121
rect 925 297 971 309
rect 925 121 931 297
rect 965 121 971 297
rect 925 109 971 121
rect 1083 297 1129 309
rect 1083 121 1089 297
rect 1123 121 1129 297
rect 1083 109 1129 121
rect 1241 297 1287 309
rect 1241 121 1247 297
rect 1281 121 1287 297
rect 1241 109 1287 121
rect 1399 297 1445 309
rect 1399 121 1405 297
rect 1439 121 1445 297
rect 1399 109 1445 121
rect 1557 297 1603 309
rect 1557 121 1563 297
rect 1597 121 1603 297
rect 1557 109 1603 121
rect 1715 297 1761 309
rect 1715 121 1721 297
rect 1755 121 1761 297
rect 1715 109 1761 121
rect 1873 297 1919 309
rect 1873 121 1879 297
rect 1913 121 1919 297
rect 1873 109 1919 121
rect 2031 297 2077 309
rect 2031 121 2037 297
rect 2071 121 2077 297
rect 2031 109 2077 121
rect 2189 297 2235 309
rect 2189 121 2195 297
rect 2229 121 2235 297
rect 2189 109 2235 121
rect 2347 297 2393 309
rect 2347 121 2353 297
rect 2387 121 2393 297
rect 2347 109 2393 121
rect -2337 71 -2245 77
rect -2337 37 -2325 71
rect -2257 37 -2245 71
rect -2337 31 -2245 37
rect -2179 71 -2087 77
rect -2179 37 -2167 71
rect -2099 37 -2087 71
rect -2179 31 -2087 37
rect -2021 71 -1929 77
rect -2021 37 -2009 71
rect -1941 37 -1929 71
rect -2021 31 -1929 37
rect -1863 71 -1771 77
rect -1863 37 -1851 71
rect -1783 37 -1771 71
rect -1863 31 -1771 37
rect -1705 71 -1613 77
rect -1705 37 -1693 71
rect -1625 37 -1613 71
rect -1705 31 -1613 37
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect 1613 71 1705 77
rect 1613 37 1625 71
rect 1693 37 1705 71
rect 1613 31 1705 37
rect 1771 71 1863 77
rect 1771 37 1783 71
rect 1851 37 1863 71
rect 1771 31 1863 37
rect 1929 71 2021 77
rect 1929 37 1941 71
rect 2009 37 2021 71
rect 1929 31 2021 37
rect 2087 71 2179 77
rect 2087 37 2099 71
rect 2167 37 2179 71
rect 2087 31 2179 37
rect 2245 71 2337 77
rect 2245 37 2257 71
rect 2325 37 2337 71
rect 2245 31 2337 37
rect -2337 -37 -2245 -31
rect -2337 -71 -2325 -37
rect -2257 -71 -2245 -37
rect -2337 -77 -2245 -71
rect -2179 -37 -2087 -31
rect -2179 -71 -2167 -37
rect -2099 -71 -2087 -37
rect -2179 -77 -2087 -71
rect -2021 -37 -1929 -31
rect -2021 -71 -2009 -37
rect -1941 -71 -1929 -37
rect -2021 -77 -1929 -71
rect -1863 -37 -1771 -31
rect -1863 -71 -1851 -37
rect -1783 -71 -1771 -37
rect -1863 -77 -1771 -71
rect -1705 -37 -1613 -31
rect -1705 -71 -1693 -37
rect -1625 -71 -1613 -37
rect -1705 -77 -1613 -71
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect 1613 -37 1705 -31
rect 1613 -71 1625 -37
rect 1693 -71 1705 -37
rect 1613 -77 1705 -71
rect 1771 -37 1863 -31
rect 1771 -71 1783 -37
rect 1851 -71 1863 -37
rect 1771 -77 1863 -71
rect 1929 -37 2021 -31
rect 1929 -71 1941 -37
rect 2009 -71 2021 -37
rect 1929 -77 2021 -71
rect 2087 -37 2179 -31
rect 2087 -71 2099 -37
rect 2167 -71 2179 -37
rect 2087 -77 2179 -71
rect 2245 -37 2337 -31
rect 2245 -71 2257 -37
rect 2325 -71 2337 -37
rect 2245 -77 2337 -71
rect -2393 -121 -2347 -109
rect -2393 -297 -2387 -121
rect -2353 -297 -2347 -121
rect -2393 -309 -2347 -297
rect -2235 -121 -2189 -109
rect -2235 -297 -2229 -121
rect -2195 -297 -2189 -121
rect -2235 -309 -2189 -297
rect -2077 -121 -2031 -109
rect -2077 -297 -2071 -121
rect -2037 -297 -2031 -121
rect -2077 -309 -2031 -297
rect -1919 -121 -1873 -109
rect -1919 -297 -1913 -121
rect -1879 -297 -1873 -121
rect -1919 -309 -1873 -297
rect -1761 -121 -1715 -109
rect -1761 -297 -1755 -121
rect -1721 -297 -1715 -121
rect -1761 -309 -1715 -297
rect -1603 -121 -1557 -109
rect -1603 -297 -1597 -121
rect -1563 -297 -1557 -121
rect -1603 -309 -1557 -297
rect -1445 -121 -1399 -109
rect -1445 -297 -1439 -121
rect -1405 -297 -1399 -121
rect -1445 -309 -1399 -297
rect -1287 -121 -1241 -109
rect -1287 -297 -1281 -121
rect -1247 -297 -1241 -121
rect -1287 -309 -1241 -297
rect -1129 -121 -1083 -109
rect -1129 -297 -1123 -121
rect -1089 -297 -1083 -121
rect -1129 -309 -1083 -297
rect -971 -121 -925 -109
rect -971 -297 -965 -121
rect -931 -297 -925 -121
rect -971 -309 -925 -297
rect -813 -121 -767 -109
rect -813 -297 -807 -121
rect -773 -297 -767 -121
rect -813 -309 -767 -297
rect -655 -121 -609 -109
rect -655 -297 -649 -121
rect -615 -297 -609 -121
rect -655 -309 -609 -297
rect -497 -121 -451 -109
rect -497 -297 -491 -121
rect -457 -297 -451 -121
rect -497 -309 -451 -297
rect -339 -121 -293 -109
rect -339 -297 -333 -121
rect -299 -297 -293 -121
rect -339 -309 -293 -297
rect -181 -121 -135 -109
rect -181 -297 -175 -121
rect -141 -297 -135 -121
rect -181 -309 -135 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 135 -121 181 -109
rect 135 -297 141 -121
rect 175 -297 181 -121
rect 135 -309 181 -297
rect 293 -121 339 -109
rect 293 -297 299 -121
rect 333 -297 339 -121
rect 293 -309 339 -297
rect 451 -121 497 -109
rect 451 -297 457 -121
rect 491 -297 497 -121
rect 451 -309 497 -297
rect 609 -121 655 -109
rect 609 -297 615 -121
rect 649 -297 655 -121
rect 609 -309 655 -297
rect 767 -121 813 -109
rect 767 -297 773 -121
rect 807 -297 813 -121
rect 767 -309 813 -297
rect 925 -121 971 -109
rect 925 -297 931 -121
rect 965 -297 971 -121
rect 925 -309 971 -297
rect 1083 -121 1129 -109
rect 1083 -297 1089 -121
rect 1123 -297 1129 -121
rect 1083 -309 1129 -297
rect 1241 -121 1287 -109
rect 1241 -297 1247 -121
rect 1281 -297 1287 -121
rect 1241 -309 1287 -297
rect 1399 -121 1445 -109
rect 1399 -297 1405 -121
rect 1439 -297 1445 -121
rect 1399 -309 1445 -297
rect 1557 -121 1603 -109
rect 1557 -297 1563 -121
rect 1597 -297 1603 -121
rect 1557 -309 1603 -297
rect 1715 -121 1761 -109
rect 1715 -297 1721 -121
rect 1755 -297 1761 -121
rect 1715 -309 1761 -297
rect 1873 -121 1919 -109
rect 1873 -297 1879 -121
rect 1913 -297 1919 -121
rect 1873 -309 1919 -297
rect 2031 -121 2077 -109
rect 2031 -297 2037 -121
rect 2071 -297 2077 -121
rect 2031 -309 2077 -297
rect 2189 -121 2235 -109
rect 2189 -297 2195 -121
rect 2229 -297 2235 -121
rect 2189 -309 2235 -297
rect 2347 -121 2393 -109
rect 2347 -297 2353 -121
rect 2387 -297 2393 -121
rect 2347 -309 2393 -297
rect -2337 -347 -2245 -341
rect -2337 -381 -2325 -347
rect -2257 -381 -2245 -347
rect -2337 -387 -2245 -381
rect -2179 -347 -2087 -341
rect -2179 -381 -2167 -347
rect -2099 -381 -2087 -347
rect -2179 -387 -2087 -381
rect -2021 -347 -1929 -341
rect -2021 -381 -2009 -347
rect -1941 -381 -1929 -347
rect -2021 -387 -1929 -381
rect -1863 -347 -1771 -341
rect -1863 -381 -1851 -347
rect -1783 -381 -1771 -347
rect -1863 -387 -1771 -381
rect -1705 -347 -1613 -341
rect -1705 -381 -1693 -347
rect -1625 -381 -1613 -347
rect -1705 -387 -1613 -381
rect -1547 -347 -1455 -341
rect -1547 -381 -1535 -347
rect -1467 -381 -1455 -347
rect -1547 -387 -1455 -381
rect -1389 -347 -1297 -341
rect -1389 -381 -1377 -347
rect -1309 -381 -1297 -347
rect -1389 -387 -1297 -381
rect -1231 -347 -1139 -341
rect -1231 -381 -1219 -347
rect -1151 -381 -1139 -347
rect -1231 -387 -1139 -381
rect -1073 -347 -981 -341
rect -1073 -381 -1061 -347
rect -993 -381 -981 -347
rect -1073 -387 -981 -381
rect -915 -347 -823 -341
rect -915 -381 -903 -347
rect -835 -381 -823 -347
rect -915 -387 -823 -381
rect -757 -347 -665 -341
rect -757 -381 -745 -347
rect -677 -381 -665 -347
rect -757 -387 -665 -381
rect -599 -347 -507 -341
rect -599 -381 -587 -347
rect -519 -381 -507 -347
rect -599 -387 -507 -381
rect -441 -347 -349 -341
rect -441 -381 -429 -347
rect -361 -381 -349 -347
rect -441 -387 -349 -381
rect -283 -347 -191 -341
rect -283 -381 -271 -347
rect -203 -381 -191 -347
rect -283 -387 -191 -381
rect -125 -347 -33 -341
rect -125 -381 -113 -347
rect -45 -381 -33 -347
rect -125 -387 -33 -381
rect 33 -347 125 -341
rect 33 -381 45 -347
rect 113 -381 125 -347
rect 33 -387 125 -381
rect 191 -347 283 -341
rect 191 -381 203 -347
rect 271 -381 283 -347
rect 191 -387 283 -381
rect 349 -347 441 -341
rect 349 -381 361 -347
rect 429 -381 441 -347
rect 349 -387 441 -381
rect 507 -347 599 -341
rect 507 -381 519 -347
rect 587 -381 599 -347
rect 507 -387 599 -381
rect 665 -347 757 -341
rect 665 -381 677 -347
rect 745 -381 757 -347
rect 665 -387 757 -381
rect 823 -347 915 -341
rect 823 -381 835 -347
rect 903 -381 915 -347
rect 823 -387 915 -381
rect 981 -347 1073 -341
rect 981 -381 993 -347
rect 1061 -381 1073 -347
rect 981 -387 1073 -381
rect 1139 -347 1231 -341
rect 1139 -381 1151 -347
rect 1219 -381 1231 -347
rect 1139 -387 1231 -381
rect 1297 -347 1389 -341
rect 1297 -381 1309 -347
rect 1377 -381 1389 -347
rect 1297 -387 1389 -381
rect 1455 -347 1547 -341
rect 1455 -381 1467 -347
rect 1535 -381 1547 -347
rect 1455 -387 1547 -381
rect 1613 -347 1705 -341
rect 1613 -381 1625 -347
rect 1693 -381 1705 -347
rect 1613 -387 1705 -381
rect 1771 -347 1863 -341
rect 1771 -381 1783 -347
rect 1851 -381 1863 -347
rect 1771 -387 1863 -381
rect 1929 -347 2021 -341
rect 1929 -381 1941 -347
rect 2009 -381 2021 -347
rect 1929 -387 2021 -381
rect 2087 -347 2179 -341
rect 2087 -381 2099 -347
rect 2167 -381 2179 -347
rect 2087 -387 2179 -381
rect 2245 -347 2337 -341
rect 2245 -381 2257 -347
rect 2325 -381 2337 -347
rect 2245 -387 2337 -381
rect -2337 -455 -2245 -449
rect -2337 -489 -2325 -455
rect -2257 -489 -2245 -455
rect -2337 -495 -2245 -489
rect -2179 -455 -2087 -449
rect -2179 -489 -2167 -455
rect -2099 -489 -2087 -455
rect -2179 -495 -2087 -489
rect -2021 -455 -1929 -449
rect -2021 -489 -2009 -455
rect -1941 -489 -1929 -455
rect -2021 -495 -1929 -489
rect -1863 -455 -1771 -449
rect -1863 -489 -1851 -455
rect -1783 -489 -1771 -455
rect -1863 -495 -1771 -489
rect -1705 -455 -1613 -449
rect -1705 -489 -1693 -455
rect -1625 -489 -1613 -455
rect -1705 -495 -1613 -489
rect -1547 -455 -1455 -449
rect -1547 -489 -1535 -455
rect -1467 -489 -1455 -455
rect -1547 -495 -1455 -489
rect -1389 -455 -1297 -449
rect -1389 -489 -1377 -455
rect -1309 -489 -1297 -455
rect -1389 -495 -1297 -489
rect -1231 -455 -1139 -449
rect -1231 -489 -1219 -455
rect -1151 -489 -1139 -455
rect -1231 -495 -1139 -489
rect -1073 -455 -981 -449
rect -1073 -489 -1061 -455
rect -993 -489 -981 -455
rect -1073 -495 -981 -489
rect -915 -455 -823 -449
rect -915 -489 -903 -455
rect -835 -489 -823 -455
rect -915 -495 -823 -489
rect -757 -455 -665 -449
rect -757 -489 -745 -455
rect -677 -489 -665 -455
rect -757 -495 -665 -489
rect -599 -455 -507 -449
rect -599 -489 -587 -455
rect -519 -489 -507 -455
rect -599 -495 -507 -489
rect -441 -455 -349 -449
rect -441 -489 -429 -455
rect -361 -489 -349 -455
rect -441 -495 -349 -489
rect -283 -455 -191 -449
rect -283 -489 -271 -455
rect -203 -489 -191 -455
rect -283 -495 -191 -489
rect -125 -455 -33 -449
rect -125 -489 -113 -455
rect -45 -489 -33 -455
rect -125 -495 -33 -489
rect 33 -455 125 -449
rect 33 -489 45 -455
rect 113 -489 125 -455
rect 33 -495 125 -489
rect 191 -455 283 -449
rect 191 -489 203 -455
rect 271 -489 283 -455
rect 191 -495 283 -489
rect 349 -455 441 -449
rect 349 -489 361 -455
rect 429 -489 441 -455
rect 349 -495 441 -489
rect 507 -455 599 -449
rect 507 -489 519 -455
rect 587 -489 599 -455
rect 507 -495 599 -489
rect 665 -455 757 -449
rect 665 -489 677 -455
rect 745 -489 757 -455
rect 665 -495 757 -489
rect 823 -455 915 -449
rect 823 -489 835 -455
rect 903 -489 915 -455
rect 823 -495 915 -489
rect 981 -455 1073 -449
rect 981 -489 993 -455
rect 1061 -489 1073 -455
rect 981 -495 1073 -489
rect 1139 -455 1231 -449
rect 1139 -489 1151 -455
rect 1219 -489 1231 -455
rect 1139 -495 1231 -489
rect 1297 -455 1389 -449
rect 1297 -489 1309 -455
rect 1377 -489 1389 -455
rect 1297 -495 1389 -489
rect 1455 -455 1547 -449
rect 1455 -489 1467 -455
rect 1535 -489 1547 -455
rect 1455 -495 1547 -489
rect 1613 -455 1705 -449
rect 1613 -489 1625 -455
rect 1693 -489 1705 -455
rect 1613 -495 1705 -489
rect 1771 -455 1863 -449
rect 1771 -489 1783 -455
rect 1851 -489 1863 -455
rect 1771 -495 1863 -489
rect 1929 -455 2021 -449
rect 1929 -489 1941 -455
rect 2009 -489 2021 -455
rect 1929 -495 2021 -489
rect 2087 -455 2179 -449
rect 2087 -489 2099 -455
rect 2167 -489 2179 -455
rect 2087 -495 2179 -489
rect 2245 -455 2337 -449
rect 2245 -489 2257 -455
rect 2325 -489 2337 -455
rect 2245 -495 2337 -489
rect -2393 -539 -2347 -527
rect -2393 -715 -2387 -539
rect -2353 -715 -2347 -539
rect -2393 -727 -2347 -715
rect -2235 -539 -2189 -527
rect -2235 -715 -2229 -539
rect -2195 -715 -2189 -539
rect -2235 -727 -2189 -715
rect -2077 -539 -2031 -527
rect -2077 -715 -2071 -539
rect -2037 -715 -2031 -539
rect -2077 -727 -2031 -715
rect -1919 -539 -1873 -527
rect -1919 -715 -1913 -539
rect -1879 -715 -1873 -539
rect -1919 -727 -1873 -715
rect -1761 -539 -1715 -527
rect -1761 -715 -1755 -539
rect -1721 -715 -1715 -539
rect -1761 -727 -1715 -715
rect -1603 -539 -1557 -527
rect -1603 -715 -1597 -539
rect -1563 -715 -1557 -539
rect -1603 -727 -1557 -715
rect -1445 -539 -1399 -527
rect -1445 -715 -1439 -539
rect -1405 -715 -1399 -539
rect -1445 -727 -1399 -715
rect -1287 -539 -1241 -527
rect -1287 -715 -1281 -539
rect -1247 -715 -1241 -539
rect -1287 -727 -1241 -715
rect -1129 -539 -1083 -527
rect -1129 -715 -1123 -539
rect -1089 -715 -1083 -539
rect -1129 -727 -1083 -715
rect -971 -539 -925 -527
rect -971 -715 -965 -539
rect -931 -715 -925 -539
rect -971 -727 -925 -715
rect -813 -539 -767 -527
rect -813 -715 -807 -539
rect -773 -715 -767 -539
rect -813 -727 -767 -715
rect -655 -539 -609 -527
rect -655 -715 -649 -539
rect -615 -715 -609 -539
rect -655 -727 -609 -715
rect -497 -539 -451 -527
rect -497 -715 -491 -539
rect -457 -715 -451 -539
rect -497 -727 -451 -715
rect -339 -539 -293 -527
rect -339 -715 -333 -539
rect -299 -715 -293 -539
rect -339 -727 -293 -715
rect -181 -539 -135 -527
rect -181 -715 -175 -539
rect -141 -715 -135 -539
rect -181 -727 -135 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 135 -539 181 -527
rect 135 -715 141 -539
rect 175 -715 181 -539
rect 135 -727 181 -715
rect 293 -539 339 -527
rect 293 -715 299 -539
rect 333 -715 339 -539
rect 293 -727 339 -715
rect 451 -539 497 -527
rect 451 -715 457 -539
rect 491 -715 497 -539
rect 451 -727 497 -715
rect 609 -539 655 -527
rect 609 -715 615 -539
rect 649 -715 655 -539
rect 609 -727 655 -715
rect 767 -539 813 -527
rect 767 -715 773 -539
rect 807 -715 813 -539
rect 767 -727 813 -715
rect 925 -539 971 -527
rect 925 -715 931 -539
rect 965 -715 971 -539
rect 925 -727 971 -715
rect 1083 -539 1129 -527
rect 1083 -715 1089 -539
rect 1123 -715 1129 -539
rect 1083 -727 1129 -715
rect 1241 -539 1287 -527
rect 1241 -715 1247 -539
rect 1281 -715 1287 -539
rect 1241 -727 1287 -715
rect 1399 -539 1445 -527
rect 1399 -715 1405 -539
rect 1439 -715 1445 -539
rect 1399 -727 1445 -715
rect 1557 -539 1603 -527
rect 1557 -715 1563 -539
rect 1597 -715 1603 -539
rect 1557 -727 1603 -715
rect 1715 -539 1761 -527
rect 1715 -715 1721 -539
rect 1755 -715 1761 -539
rect 1715 -727 1761 -715
rect 1873 -539 1919 -527
rect 1873 -715 1879 -539
rect 1913 -715 1919 -539
rect 1873 -727 1919 -715
rect 2031 -539 2077 -527
rect 2031 -715 2037 -539
rect 2071 -715 2077 -539
rect 2031 -727 2077 -715
rect 2189 -539 2235 -527
rect 2189 -715 2195 -539
rect 2229 -715 2235 -539
rect 2189 -727 2235 -715
rect 2347 -539 2393 -527
rect 2347 -715 2353 -539
rect 2387 -715 2393 -539
rect 2347 -727 2393 -715
rect -2337 -765 -2245 -759
rect -2337 -799 -2325 -765
rect -2257 -799 -2245 -765
rect -2337 -805 -2245 -799
rect -2179 -765 -2087 -759
rect -2179 -799 -2167 -765
rect -2099 -799 -2087 -765
rect -2179 -805 -2087 -799
rect -2021 -765 -1929 -759
rect -2021 -799 -2009 -765
rect -1941 -799 -1929 -765
rect -2021 -805 -1929 -799
rect -1863 -765 -1771 -759
rect -1863 -799 -1851 -765
rect -1783 -799 -1771 -765
rect -1863 -805 -1771 -799
rect -1705 -765 -1613 -759
rect -1705 -799 -1693 -765
rect -1625 -799 -1613 -765
rect -1705 -805 -1613 -799
rect -1547 -765 -1455 -759
rect -1547 -799 -1535 -765
rect -1467 -799 -1455 -765
rect -1547 -805 -1455 -799
rect -1389 -765 -1297 -759
rect -1389 -799 -1377 -765
rect -1309 -799 -1297 -765
rect -1389 -805 -1297 -799
rect -1231 -765 -1139 -759
rect -1231 -799 -1219 -765
rect -1151 -799 -1139 -765
rect -1231 -805 -1139 -799
rect -1073 -765 -981 -759
rect -1073 -799 -1061 -765
rect -993 -799 -981 -765
rect -1073 -805 -981 -799
rect -915 -765 -823 -759
rect -915 -799 -903 -765
rect -835 -799 -823 -765
rect -915 -805 -823 -799
rect -757 -765 -665 -759
rect -757 -799 -745 -765
rect -677 -799 -665 -765
rect -757 -805 -665 -799
rect -599 -765 -507 -759
rect -599 -799 -587 -765
rect -519 -799 -507 -765
rect -599 -805 -507 -799
rect -441 -765 -349 -759
rect -441 -799 -429 -765
rect -361 -799 -349 -765
rect -441 -805 -349 -799
rect -283 -765 -191 -759
rect -283 -799 -271 -765
rect -203 -799 -191 -765
rect -283 -805 -191 -799
rect -125 -765 -33 -759
rect -125 -799 -113 -765
rect -45 -799 -33 -765
rect -125 -805 -33 -799
rect 33 -765 125 -759
rect 33 -799 45 -765
rect 113 -799 125 -765
rect 33 -805 125 -799
rect 191 -765 283 -759
rect 191 -799 203 -765
rect 271 -799 283 -765
rect 191 -805 283 -799
rect 349 -765 441 -759
rect 349 -799 361 -765
rect 429 -799 441 -765
rect 349 -805 441 -799
rect 507 -765 599 -759
rect 507 -799 519 -765
rect 587 -799 599 -765
rect 507 -805 599 -799
rect 665 -765 757 -759
rect 665 -799 677 -765
rect 745 -799 757 -765
rect 665 -805 757 -799
rect 823 -765 915 -759
rect 823 -799 835 -765
rect 903 -799 915 -765
rect 823 -805 915 -799
rect 981 -765 1073 -759
rect 981 -799 993 -765
rect 1061 -799 1073 -765
rect 981 -805 1073 -799
rect 1139 -765 1231 -759
rect 1139 -799 1151 -765
rect 1219 -799 1231 -765
rect 1139 -805 1231 -799
rect 1297 -765 1389 -759
rect 1297 -799 1309 -765
rect 1377 -799 1389 -765
rect 1297 -805 1389 -799
rect 1455 -765 1547 -759
rect 1455 -799 1467 -765
rect 1535 -799 1547 -765
rect 1455 -805 1547 -799
rect 1613 -765 1705 -759
rect 1613 -799 1625 -765
rect 1693 -799 1705 -765
rect 1613 -805 1705 -799
rect 1771 -765 1863 -759
rect 1771 -799 1783 -765
rect 1851 -799 1863 -765
rect 1771 -805 1863 -799
rect 1929 -765 2021 -759
rect 1929 -799 1941 -765
rect 2009 -799 2021 -765
rect 1929 -805 2021 -799
rect 2087 -765 2179 -759
rect 2087 -799 2099 -765
rect 2167 -799 2179 -765
rect 2087 -805 2179 -799
rect 2245 -765 2337 -759
rect 2245 -799 2257 -765
rect 2325 -799 2337 -765
rect 2245 -805 2337 -799
<< properties >>
string FIXED_BBOX -2504 -920 2504 920
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 4 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
