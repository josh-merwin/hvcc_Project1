magic
tech sky130B
magscale 1 2
timestamp 1651944383
<< nwell >>
rect -16029 -397 16029 397
<< mvpmos >>
rect -15771 -100 -15671 100
rect -15613 -100 -15513 100
rect -15455 -100 -15355 100
rect -15297 -100 -15197 100
rect -15139 -100 -15039 100
rect -14981 -100 -14881 100
rect -14823 -100 -14723 100
rect -14665 -100 -14565 100
rect -14507 -100 -14407 100
rect -14349 -100 -14249 100
rect -14191 -100 -14091 100
rect -14033 -100 -13933 100
rect -13875 -100 -13775 100
rect -13717 -100 -13617 100
rect -13559 -100 -13459 100
rect -13401 -100 -13301 100
rect -13243 -100 -13143 100
rect -13085 -100 -12985 100
rect -12927 -100 -12827 100
rect -12769 -100 -12669 100
rect -12611 -100 -12511 100
rect -12453 -100 -12353 100
rect -12295 -100 -12195 100
rect -12137 -100 -12037 100
rect -11979 -100 -11879 100
rect -11821 -100 -11721 100
rect -11663 -100 -11563 100
rect -11505 -100 -11405 100
rect -11347 -100 -11247 100
rect -11189 -100 -11089 100
rect -11031 -100 -10931 100
rect -10873 -100 -10773 100
rect -10715 -100 -10615 100
rect -10557 -100 -10457 100
rect -10399 -100 -10299 100
rect -10241 -100 -10141 100
rect -10083 -100 -9983 100
rect -9925 -100 -9825 100
rect -9767 -100 -9667 100
rect -9609 -100 -9509 100
rect -9451 -100 -9351 100
rect -9293 -100 -9193 100
rect -9135 -100 -9035 100
rect -8977 -100 -8877 100
rect -8819 -100 -8719 100
rect -8661 -100 -8561 100
rect -8503 -100 -8403 100
rect -8345 -100 -8245 100
rect -8187 -100 -8087 100
rect -8029 -100 -7929 100
rect -7871 -100 -7771 100
rect -7713 -100 -7613 100
rect -7555 -100 -7455 100
rect -7397 -100 -7297 100
rect -7239 -100 -7139 100
rect -7081 -100 -6981 100
rect -6923 -100 -6823 100
rect -6765 -100 -6665 100
rect -6607 -100 -6507 100
rect -6449 -100 -6349 100
rect -6291 -100 -6191 100
rect -6133 -100 -6033 100
rect -5975 -100 -5875 100
rect -5817 -100 -5717 100
rect -5659 -100 -5559 100
rect -5501 -100 -5401 100
rect -5343 -100 -5243 100
rect -5185 -100 -5085 100
rect -5027 -100 -4927 100
rect -4869 -100 -4769 100
rect -4711 -100 -4611 100
rect -4553 -100 -4453 100
rect -4395 -100 -4295 100
rect -4237 -100 -4137 100
rect -4079 -100 -3979 100
rect -3921 -100 -3821 100
rect -3763 -100 -3663 100
rect -3605 -100 -3505 100
rect -3447 -100 -3347 100
rect -3289 -100 -3189 100
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect 3189 -100 3289 100
rect 3347 -100 3447 100
rect 3505 -100 3605 100
rect 3663 -100 3763 100
rect 3821 -100 3921 100
rect 3979 -100 4079 100
rect 4137 -100 4237 100
rect 4295 -100 4395 100
rect 4453 -100 4553 100
rect 4611 -100 4711 100
rect 4769 -100 4869 100
rect 4927 -100 5027 100
rect 5085 -100 5185 100
rect 5243 -100 5343 100
rect 5401 -100 5501 100
rect 5559 -100 5659 100
rect 5717 -100 5817 100
rect 5875 -100 5975 100
rect 6033 -100 6133 100
rect 6191 -100 6291 100
rect 6349 -100 6449 100
rect 6507 -100 6607 100
rect 6665 -100 6765 100
rect 6823 -100 6923 100
rect 6981 -100 7081 100
rect 7139 -100 7239 100
rect 7297 -100 7397 100
rect 7455 -100 7555 100
rect 7613 -100 7713 100
rect 7771 -100 7871 100
rect 7929 -100 8029 100
rect 8087 -100 8187 100
rect 8245 -100 8345 100
rect 8403 -100 8503 100
rect 8561 -100 8661 100
rect 8719 -100 8819 100
rect 8877 -100 8977 100
rect 9035 -100 9135 100
rect 9193 -100 9293 100
rect 9351 -100 9451 100
rect 9509 -100 9609 100
rect 9667 -100 9767 100
rect 9825 -100 9925 100
rect 9983 -100 10083 100
rect 10141 -100 10241 100
rect 10299 -100 10399 100
rect 10457 -100 10557 100
rect 10615 -100 10715 100
rect 10773 -100 10873 100
rect 10931 -100 11031 100
rect 11089 -100 11189 100
rect 11247 -100 11347 100
rect 11405 -100 11505 100
rect 11563 -100 11663 100
rect 11721 -100 11821 100
rect 11879 -100 11979 100
rect 12037 -100 12137 100
rect 12195 -100 12295 100
rect 12353 -100 12453 100
rect 12511 -100 12611 100
rect 12669 -100 12769 100
rect 12827 -100 12927 100
rect 12985 -100 13085 100
rect 13143 -100 13243 100
rect 13301 -100 13401 100
rect 13459 -100 13559 100
rect 13617 -100 13717 100
rect 13775 -100 13875 100
rect 13933 -100 14033 100
rect 14091 -100 14191 100
rect 14249 -100 14349 100
rect 14407 -100 14507 100
rect 14565 -100 14665 100
rect 14723 -100 14823 100
rect 14881 -100 14981 100
rect 15039 -100 15139 100
rect 15197 -100 15297 100
rect 15355 -100 15455 100
rect 15513 -100 15613 100
rect 15671 -100 15771 100
<< mvpdiff >>
rect -15829 88 -15771 100
rect -15829 -88 -15817 88
rect -15783 -88 -15771 88
rect -15829 -100 -15771 -88
rect -15671 88 -15613 100
rect -15671 -88 -15659 88
rect -15625 -88 -15613 88
rect -15671 -100 -15613 -88
rect -15513 88 -15455 100
rect -15513 -88 -15501 88
rect -15467 -88 -15455 88
rect -15513 -100 -15455 -88
rect -15355 88 -15297 100
rect -15355 -88 -15343 88
rect -15309 -88 -15297 88
rect -15355 -100 -15297 -88
rect -15197 88 -15139 100
rect -15197 -88 -15185 88
rect -15151 -88 -15139 88
rect -15197 -100 -15139 -88
rect -15039 88 -14981 100
rect -15039 -88 -15027 88
rect -14993 -88 -14981 88
rect -15039 -100 -14981 -88
rect -14881 88 -14823 100
rect -14881 -88 -14869 88
rect -14835 -88 -14823 88
rect -14881 -100 -14823 -88
rect -14723 88 -14665 100
rect -14723 -88 -14711 88
rect -14677 -88 -14665 88
rect -14723 -100 -14665 -88
rect -14565 88 -14507 100
rect -14565 -88 -14553 88
rect -14519 -88 -14507 88
rect -14565 -100 -14507 -88
rect -14407 88 -14349 100
rect -14407 -88 -14395 88
rect -14361 -88 -14349 88
rect -14407 -100 -14349 -88
rect -14249 88 -14191 100
rect -14249 -88 -14237 88
rect -14203 -88 -14191 88
rect -14249 -100 -14191 -88
rect -14091 88 -14033 100
rect -14091 -88 -14079 88
rect -14045 -88 -14033 88
rect -14091 -100 -14033 -88
rect -13933 88 -13875 100
rect -13933 -88 -13921 88
rect -13887 -88 -13875 88
rect -13933 -100 -13875 -88
rect -13775 88 -13717 100
rect -13775 -88 -13763 88
rect -13729 -88 -13717 88
rect -13775 -100 -13717 -88
rect -13617 88 -13559 100
rect -13617 -88 -13605 88
rect -13571 -88 -13559 88
rect -13617 -100 -13559 -88
rect -13459 88 -13401 100
rect -13459 -88 -13447 88
rect -13413 -88 -13401 88
rect -13459 -100 -13401 -88
rect -13301 88 -13243 100
rect -13301 -88 -13289 88
rect -13255 -88 -13243 88
rect -13301 -100 -13243 -88
rect -13143 88 -13085 100
rect -13143 -88 -13131 88
rect -13097 -88 -13085 88
rect -13143 -100 -13085 -88
rect -12985 88 -12927 100
rect -12985 -88 -12973 88
rect -12939 -88 -12927 88
rect -12985 -100 -12927 -88
rect -12827 88 -12769 100
rect -12827 -88 -12815 88
rect -12781 -88 -12769 88
rect -12827 -100 -12769 -88
rect -12669 88 -12611 100
rect -12669 -88 -12657 88
rect -12623 -88 -12611 88
rect -12669 -100 -12611 -88
rect -12511 88 -12453 100
rect -12511 -88 -12499 88
rect -12465 -88 -12453 88
rect -12511 -100 -12453 -88
rect -12353 88 -12295 100
rect -12353 -88 -12341 88
rect -12307 -88 -12295 88
rect -12353 -100 -12295 -88
rect -12195 88 -12137 100
rect -12195 -88 -12183 88
rect -12149 -88 -12137 88
rect -12195 -100 -12137 -88
rect -12037 88 -11979 100
rect -12037 -88 -12025 88
rect -11991 -88 -11979 88
rect -12037 -100 -11979 -88
rect -11879 88 -11821 100
rect -11879 -88 -11867 88
rect -11833 -88 -11821 88
rect -11879 -100 -11821 -88
rect -11721 88 -11663 100
rect -11721 -88 -11709 88
rect -11675 -88 -11663 88
rect -11721 -100 -11663 -88
rect -11563 88 -11505 100
rect -11563 -88 -11551 88
rect -11517 -88 -11505 88
rect -11563 -100 -11505 -88
rect -11405 88 -11347 100
rect -11405 -88 -11393 88
rect -11359 -88 -11347 88
rect -11405 -100 -11347 -88
rect -11247 88 -11189 100
rect -11247 -88 -11235 88
rect -11201 -88 -11189 88
rect -11247 -100 -11189 -88
rect -11089 88 -11031 100
rect -11089 -88 -11077 88
rect -11043 -88 -11031 88
rect -11089 -100 -11031 -88
rect -10931 88 -10873 100
rect -10931 -88 -10919 88
rect -10885 -88 -10873 88
rect -10931 -100 -10873 -88
rect -10773 88 -10715 100
rect -10773 -88 -10761 88
rect -10727 -88 -10715 88
rect -10773 -100 -10715 -88
rect -10615 88 -10557 100
rect -10615 -88 -10603 88
rect -10569 -88 -10557 88
rect -10615 -100 -10557 -88
rect -10457 88 -10399 100
rect -10457 -88 -10445 88
rect -10411 -88 -10399 88
rect -10457 -100 -10399 -88
rect -10299 88 -10241 100
rect -10299 -88 -10287 88
rect -10253 -88 -10241 88
rect -10299 -100 -10241 -88
rect -10141 88 -10083 100
rect -10141 -88 -10129 88
rect -10095 -88 -10083 88
rect -10141 -100 -10083 -88
rect -9983 88 -9925 100
rect -9983 -88 -9971 88
rect -9937 -88 -9925 88
rect -9983 -100 -9925 -88
rect -9825 88 -9767 100
rect -9825 -88 -9813 88
rect -9779 -88 -9767 88
rect -9825 -100 -9767 -88
rect -9667 88 -9609 100
rect -9667 -88 -9655 88
rect -9621 -88 -9609 88
rect -9667 -100 -9609 -88
rect -9509 88 -9451 100
rect -9509 -88 -9497 88
rect -9463 -88 -9451 88
rect -9509 -100 -9451 -88
rect -9351 88 -9293 100
rect -9351 -88 -9339 88
rect -9305 -88 -9293 88
rect -9351 -100 -9293 -88
rect -9193 88 -9135 100
rect -9193 -88 -9181 88
rect -9147 -88 -9135 88
rect -9193 -100 -9135 -88
rect -9035 88 -8977 100
rect -9035 -88 -9023 88
rect -8989 -88 -8977 88
rect -9035 -100 -8977 -88
rect -8877 88 -8819 100
rect -8877 -88 -8865 88
rect -8831 -88 -8819 88
rect -8877 -100 -8819 -88
rect -8719 88 -8661 100
rect -8719 -88 -8707 88
rect -8673 -88 -8661 88
rect -8719 -100 -8661 -88
rect -8561 88 -8503 100
rect -8561 -88 -8549 88
rect -8515 -88 -8503 88
rect -8561 -100 -8503 -88
rect -8403 88 -8345 100
rect -8403 -88 -8391 88
rect -8357 -88 -8345 88
rect -8403 -100 -8345 -88
rect -8245 88 -8187 100
rect -8245 -88 -8233 88
rect -8199 -88 -8187 88
rect -8245 -100 -8187 -88
rect -8087 88 -8029 100
rect -8087 -88 -8075 88
rect -8041 -88 -8029 88
rect -8087 -100 -8029 -88
rect -7929 88 -7871 100
rect -7929 -88 -7917 88
rect -7883 -88 -7871 88
rect -7929 -100 -7871 -88
rect -7771 88 -7713 100
rect -7771 -88 -7759 88
rect -7725 -88 -7713 88
rect -7771 -100 -7713 -88
rect -7613 88 -7555 100
rect -7613 -88 -7601 88
rect -7567 -88 -7555 88
rect -7613 -100 -7555 -88
rect -7455 88 -7397 100
rect -7455 -88 -7443 88
rect -7409 -88 -7397 88
rect -7455 -100 -7397 -88
rect -7297 88 -7239 100
rect -7297 -88 -7285 88
rect -7251 -88 -7239 88
rect -7297 -100 -7239 -88
rect -7139 88 -7081 100
rect -7139 -88 -7127 88
rect -7093 -88 -7081 88
rect -7139 -100 -7081 -88
rect -6981 88 -6923 100
rect -6981 -88 -6969 88
rect -6935 -88 -6923 88
rect -6981 -100 -6923 -88
rect -6823 88 -6765 100
rect -6823 -88 -6811 88
rect -6777 -88 -6765 88
rect -6823 -100 -6765 -88
rect -6665 88 -6607 100
rect -6665 -88 -6653 88
rect -6619 -88 -6607 88
rect -6665 -100 -6607 -88
rect -6507 88 -6449 100
rect -6507 -88 -6495 88
rect -6461 -88 -6449 88
rect -6507 -100 -6449 -88
rect -6349 88 -6291 100
rect -6349 -88 -6337 88
rect -6303 -88 -6291 88
rect -6349 -100 -6291 -88
rect -6191 88 -6133 100
rect -6191 -88 -6179 88
rect -6145 -88 -6133 88
rect -6191 -100 -6133 -88
rect -6033 88 -5975 100
rect -6033 -88 -6021 88
rect -5987 -88 -5975 88
rect -6033 -100 -5975 -88
rect -5875 88 -5817 100
rect -5875 -88 -5863 88
rect -5829 -88 -5817 88
rect -5875 -100 -5817 -88
rect -5717 88 -5659 100
rect -5717 -88 -5705 88
rect -5671 -88 -5659 88
rect -5717 -100 -5659 -88
rect -5559 88 -5501 100
rect -5559 -88 -5547 88
rect -5513 -88 -5501 88
rect -5559 -100 -5501 -88
rect -5401 88 -5343 100
rect -5401 -88 -5389 88
rect -5355 -88 -5343 88
rect -5401 -100 -5343 -88
rect -5243 88 -5185 100
rect -5243 -88 -5231 88
rect -5197 -88 -5185 88
rect -5243 -100 -5185 -88
rect -5085 88 -5027 100
rect -5085 -88 -5073 88
rect -5039 -88 -5027 88
rect -5085 -100 -5027 -88
rect -4927 88 -4869 100
rect -4927 -88 -4915 88
rect -4881 -88 -4869 88
rect -4927 -100 -4869 -88
rect -4769 88 -4711 100
rect -4769 -88 -4757 88
rect -4723 -88 -4711 88
rect -4769 -100 -4711 -88
rect -4611 88 -4553 100
rect -4611 -88 -4599 88
rect -4565 -88 -4553 88
rect -4611 -100 -4553 -88
rect -4453 88 -4395 100
rect -4453 -88 -4441 88
rect -4407 -88 -4395 88
rect -4453 -100 -4395 -88
rect -4295 88 -4237 100
rect -4295 -88 -4283 88
rect -4249 -88 -4237 88
rect -4295 -100 -4237 -88
rect -4137 88 -4079 100
rect -4137 -88 -4125 88
rect -4091 -88 -4079 88
rect -4137 -100 -4079 -88
rect -3979 88 -3921 100
rect -3979 -88 -3967 88
rect -3933 -88 -3921 88
rect -3979 -100 -3921 -88
rect -3821 88 -3763 100
rect -3821 -88 -3809 88
rect -3775 -88 -3763 88
rect -3821 -100 -3763 -88
rect -3663 88 -3605 100
rect -3663 -88 -3651 88
rect -3617 -88 -3605 88
rect -3663 -100 -3605 -88
rect -3505 88 -3447 100
rect -3505 -88 -3493 88
rect -3459 -88 -3447 88
rect -3505 -100 -3447 -88
rect -3347 88 -3289 100
rect -3347 -88 -3335 88
rect -3301 -88 -3289 88
rect -3347 -100 -3289 -88
rect -3189 88 -3131 100
rect -3189 -88 -3177 88
rect -3143 -88 -3131 88
rect -3189 -100 -3131 -88
rect -3031 88 -2973 100
rect -3031 -88 -3019 88
rect -2985 -88 -2973 88
rect -3031 -100 -2973 -88
rect -2873 88 -2815 100
rect -2873 -88 -2861 88
rect -2827 -88 -2815 88
rect -2873 -100 -2815 -88
rect -2715 88 -2657 100
rect -2715 -88 -2703 88
rect -2669 -88 -2657 88
rect -2715 -100 -2657 -88
rect -2557 88 -2499 100
rect -2557 -88 -2545 88
rect -2511 -88 -2499 88
rect -2557 -100 -2499 -88
rect -2399 88 -2341 100
rect -2399 -88 -2387 88
rect -2353 -88 -2341 88
rect -2399 -100 -2341 -88
rect -2241 88 -2183 100
rect -2241 -88 -2229 88
rect -2195 -88 -2183 88
rect -2241 -100 -2183 -88
rect -2083 88 -2025 100
rect -2083 -88 -2071 88
rect -2037 -88 -2025 88
rect -2083 -100 -2025 -88
rect -1925 88 -1867 100
rect -1925 -88 -1913 88
rect -1879 -88 -1867 88
rect -1925 -100 -1867 -88
rect -1767 88 -1709 100
rect -1767 -88 -1755 88
rect -1721 -88 -1709 88
rect -1767 -100 -1709 -88
rect -1609 88 -1551 100
rect -1609 -88 -1597 88
rect -1563 -88 -1551 88
rect -1609 -100 -1551 -88
rect -1451 88 -1393 100
rect -1451 -88 -1439 88
rect -1405 -88 -1393 88
rect -1451 -100 -1393 -88
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
rect 1393 88 1451 100
rect 1393 -88 1405 88
rect 1439 -88 1451 88
rect 1393 -100 1451 -88
rect 1551 88 1609 100
rect 1551 -88 1563 88
rect 1597 -88 1609 88
rect 1551 -100 1609 -88
rect 1709 88 1767 100
rect 1709 -88 1721 88
rect 1755 -88 1767 88
rect 1709 -100 1767 -88
rect 1867 88 1925 100
rect 1867 -88 1879 88
rect 1913 -88 1925 88
rect 1867 -100 1925 -88
rect 2025 88 2083 100
rect 2025 -88 2037 88
rect 2071 -88 2083 88
rect 2025 -100 2083 -88
rect 2183 88 2241 100
rect 2183 -88 2195 88
rect 2229 -88 2241 88
rect 2183 -100 2241 -88
rect 2341 88 2399 100
rect 2341 -88 2353 88
rect 2387 -88 2399 88
rect 2341 -100 2399 -88
rect 2499 88 2557 100
rect 2499 -88 2511 88
rect 2545 -88 2557 88
rect 2499 -100 2557 -88
rect 2657 88 2715 100
rect 2657 -88 2669 88
rect 2703 -88 2715 88
rect 2657 -100 2715 -88
rect 2815 88 2873 100
rect 2815 -88 2827 88
rect 2861 -88 2873 88
rect 2815 -100 2873 -88
rect 2973 88 3031 100
rect 2973 -88 2985 88
rect 3019 -88 3031 88
rect 2973 -100 3031 -88
rect 3131 88 3189 100
rect 3131 -88 3143 88
rect 3177 -88 3189 88
rect 3131 -100 3189 -88
rect 3289 88 3347 100
rect 3289 -88 3301 88
rect 3335 -88 3347 88
rect 3289 -100 3347 -88
rect 3447 88 3505 100
rect 3447 -88 3459 88
rect 3493 -88 3505 88
rect 3447 -100 3505 -88
rect 3605 88 3663 100
rect 3605 -88 3617 88
rect 3651 -88 3663 88
rect 3605 -100 3663 -88
rect 3763 88 3821 100
rect 3763 -88 3775 88
rect 3809 -88 3821 88
rect 3763 -100 3821 -88
rect 3921 88 3979 100
rect 3921 -88 3933 88
rect 3967 -88 3979 88
rect 3921 -100 3979 -88
rect 4079 88 4137 100
rect 4079 -88 4091 88
rect 4125 -88 4137 88
rect 4079 -100 4137 -88
rect 4237 88 4295 100
rect 4237 -88 4249 88
rect 4283 -88 4295 88
rect 4237 -100 4295 -88
rect 4395 88 4453 100
rect 4395 -88 4407 88
rect 4441 -88 4453 88
rect 4395 -100 4453 -88
rect 4553 88 4611 100
rect 4553 -88 4565 88
rect 4599 -88 4611 88
rect 4553 -100 4611 -88
rect 4711 88 4769 100
rect 4711 -88 4723 88
rect 4757 -88 4769 88
rect 4711 -100 4769 -88
rect 4869 88 4927 100
rect 4869 -88 4881 88
rect 4915 -88 4927 88
rect 4869 -100 4927 -88
rect 5027 88 5085 100
rect 5027 -88 5039 88
rect 5073 -88 5085 88
rect 5027 -100 5085 -88
rect 5185 88 5243 100
rect 5185 -88 5197 88
rect 5231 -88 5243 88
rect 5185 -100 5243 -88
rect 5343 88 5401 100
rect 5343 -88 5355 88
rect 5389 -88 5401 88
rect 5343 -100 5401 -88
rect 5501 88 5559 100
rect 5501 -88 5513 88
rect 5547 -88 5559 88
rect 5501 -100 5559 -88
rect 5659 88 5717 100
rect 5659 -88 5671 88
rect 5705 -88 5717 88
rect 5659 -100 5717 -88
rect 5817 88 5875 100
rect 5817 -88 5829 88
rect 5863 -88 5875 88
rect 5817 -100 5875 -88
rect 5975 88 6033 100
rect 5975 -88 5987 88
rect 6021 -88 6033 88
rect 5975 -100 6033 -88
rect 6133 88 6191 100
rect 6133 -88 6145 88
rect 6179 -88 6191 88
rect 6133 -100 6191 -88
rect 6291 88 6349 100
rect 6291 -88 6303 88
rect 6337 -88 6349 88
rect 6291 -100 6349 -88
rect 6449 88 6507 100
rect 6449 -88 6461 88
rect 6495 -88 6507 88
rect 6449 -100 6507 -88
rect 6607 88 6665 100
rect 6607 -88 6619 88
rect 6653 -88 6665 88
rect 6607 -100 6665 -88
rect 6765 88 6823 100
rect 6765 -88 6777 88
rect 6811 -88 6823 88
rect 6765 -100 6823 -88
rect 6923 88 6981 100
rect 6923 -88 6935 88
rect 6969 -88 6981 88
rect 6923 -100 6981 -88
rect 7081 88 7139 100
rect 7081 -88 7093 88
rect 7127 -88 7139 88
rect 7081 -100 7139 -88
rect 7239 88 7297 100
rect 7239 -88 7251 88
rect 7285 -88 7297 88
rect 7239 -100 7297 -88
rect 7397 88 7455 100
rect 7397 -88 7409 88
rect 7443 -88 7455 88
rect 7397 -100 7455 -88
rect 7555 88 7613 100
rect 7555 -88 7567 88
rect 7601 -88 7613 88
rect 7555 -100 7613 -88
rect 7713 88 7771 100
rect 7713 -88 7725 88
rect 7759 -88 7771 88
rect 7713 -100 7771 -88
rect 7871 88 7929 100
rect 7871 -88 7883 88
rect 7917 -88 7929 88
rect 7871 -100 7929 -88
rect 8029 88 8087 100
rect 8029 -88 8041 88
rect 8075 -88 8087 88
rect 8029 -100 8087 -88
rect 8187 88 8245 100
rect 8187 -88 8199 88
rect 8233 -88 8245 88
rect 8187 -100 8245 -88
rect 8345 88 8403 100
rect 8345 -88 8357 88
rect 8391 -88 8403 88
rect 8345 -100 8403 -88
rect 8503 88 8561 100
rect 8503 -88 8515 88
rect 8549 -88 8561 88
rect 8503 -100 8561 -88
rect 8661 88 8719 100
rect 8661 -88 8673 88
rect 8707 -88 8719 88
rect 8661 -100 8719 -88
rect 8819 88 8877 100
rect 8819 -88 8831 88
rect 8865 -88 8877 88
rect 8819 -100 8877 -88
rect 8977 88 9035 100
rect 8977 -88 8989 88
rect 9023 -88 9035 88
rect 8977 -100 9035 -88
rect 9135 88 9193 100
rect 9135 -88 9147 88
rect 9181 -88 9193 88
rect 9135 -100 9193 -88
rect 9293 88 9351 100
rect 9293 -88 9305 88
rect 9339 -88 9351 88
rect 9293 -100 9351 -88
rect 9451 88 9509 100
rect 9451 -88 9463 88
rect 9497 -88 9509 88
rect 9451 -100 9509 -88
rect 9609 88 9667 100
rect 9609 -88 9621 88
rect 9655 -88 9667 88
rect 9609 -100 9667 -88
rect 9767 88 9825 100
rect 9767 -88 9779 88
rect 9813 -88 9825 88
rect 9767 -100 9825 -88
rect 9925 88 9983 100
rect 9925 -88 9937 88
rect 9971 -88 9983 88
rect 9925 -100 9983 -88
rect 10083 88 10141 100
rect 10083 -88 10095 88
rect 10129 -88 10141 88
rect 10083 -100 10141 -88
rect 10241 88 10299 100
rect 10241 -88 10253 88
rect 10287 -88 10299 88
rect 10241 -100 10299 -88
rect 10399 88 10457 100
rect 10399 -88 10411 88
rect 10445 -88 10457 88
rect 10399 -100 10457 -88
rect 10557 88 10615 100
rect 10557 -88 10569 88
rect 10603 -88 10615 88
rect 10557 -100 10615 -88
rect 10715 88 10773 100
rect 10715 -88 10727 88
rect 10761 -88 10773 88
rect 10715 -100 10773 -88
rect 10873 88 10931 100
rect 10873 -88 10885 88
rect 10919 -88 10931 88
rect 10873 -100 10931 -88
rect 11031 88 11089 100
rect 11031 -88 11043 88
rect 11077 -88 11089 88
rect 11031 -100 11089 -88
rect 11189 88 11247 100
rect 11189 -88 11201 88
rect 11235 -88 11247 88
rect 11189 -100 11247 -88
rect 11347 88 11405 100
rect 11347 -88 11359 88
rect 11393 -88 11405 88
rect 11347 -100 11405 -88
rect 11505 88 11563 100
rect 11505 -88 11517 88
rect 11551 -88 11563 88
rect 11505 -100 11563 -88
rect 11663 88 11721 100
rect 11663 -88 11675 88
rect 11709 -88 11721 88
rect 11663 -100 11721 -88
rect 11821 88 11879 100
rect 11821 -88 11833 88
rect 11867 -88 11879 88
rect 11821 -100 11879 -88
rect 11979 88 12037 100
rect 11979 -88 11991 88
rect 12025 -88 12037 88
rect 11979 -100 12037 -88
rect 12137 88 12195 100
rect 12137 -88 12149 88
rect 12183 -88 12195 88
rect 12137 -100 12195 -88
rect 12295 88 12353 100
rect 12295 -88 12307 88
rect 12341 -88 12353 88
rect 12295 -100 12353 -88
rect 12453 88 12511 100
rect 12453 -88 12465 88
rect 12499 -88 12511 88
rect 12453 -100 12511 -88
rect 12611 88 12669 100
rect 12611 -88 12623 88
rect 12657 -88 12669 88
rect 12611 -100 12669 -88
rect 12769 88 12827 100
rect 12769 -88 12781 88
rect 12815 -88 12827 88
rect 12769 -100 12827 -88
rect 12927 88 12985 100
rect 12927 -88 12939 88
rect 12973 -88 12985 88
rect 12927 -100 12985 -88
rect 13085 88 13143 100
rect 13085 -88 13097 88
rect 13131 -88 13143 88
rect 13085 -100 13143 -88
rect 13243 88 13301 100
rect 13243 -88 13255 88
rect 13289 -88 13301 88
rect 13243 -100 13301 -88
rect 13401 88 13459 100
rect 13401 -88 13413 88
rect 13447 -88 13459 88
rect 13401 -100 13459 -88
rect 13559 88 13617 100
rect 13559 -88 13571 88
rect 13605 -88 13617 88
rect 13559 -100 13617 -88
rect 13717 88 13775 100
rect 13717 -88 13729 88
rect 13763 -88 13775 88
rect 13717 -100 13775 -88
rect 13875 88 13933 100
rect 13875 -88 13887 88
rect 13921 -88 13933 88
rect 13875 -100 13933 -88
rect 14033 88 14091 100
rect 14033 -88 14045 88
rect 14079 -88 14091 88
rect 14033 -100 14091 -88
rect 14191 88 14249 100
rect 14191 -88 14203 88
rect 14237 -88 14249 88
rect 14191 -100 14249 -88
rect 14349 88 14407 100
rect 14349 -88 14361 88
rect 14395 -88 14407 88
rect 14349 -100 14407 -88
rect 14507 88 14565 100
rect 14507 -88 14519 88
rect 14553 -88 14565 88
rect 14507 -100 14565 -88
rect 14665 88 14723 100
rect 14665 -88 14677 88
rect 14711 -88 14723 88
rect 14665 -100 14723 -88
rect 14823 88 14881 100
rect 14823 -88 14835 88
rect 14869 -88 14881 88
rect 14823 -100 14881 -88
rect 14981 88 15039 100
rect 14981 -88 14993 88
rect 15027 -88 15039 88
rect 14981 -100 15039 -88
rect 15139 88 15197 100
rect 15139 -88 15151 88
rect 15185 -88 15197 88
rect 15139 -100 15197 -88
rect 15297 88 15355 100
rect 15297 -88 15309 88
rect 15343 -88 15355 88
rect 15297 -100 15355 -88
rect 15455 88 15513 100
rect 15455 -88 15467 88
rect 15501 -88 15513 88
rect 15455 -100 15513 -88
rect 15613 88 15671 100
rect 15613 -88 15625 88
rect 15659 -88 15671 88
rect 15613 -100 15671 -88
rect 15771 88 15829 100
rect 15771 -88 15783 88
rect 15817 -88 15829 88
rect 15771 -100 15829 -88
<< mvpdiffc >>
rect -15817 -88 -15783 88
rect -15659 -88 -15625 88
rect -15501 -88 -15467 88
rect -15343 -88 -15309 88
rect -15185 -88 -15151 88
rect -15027 -88 -14993 88
rect -14869 -88 -14835 88
rect -14711 -88 -14677 88
rect -14553 -88 -14519 88
rect -14395 -88 -14361 88
rect -14237 -88 -14203 88
rect -14079 -88 -14045 88
rect -13921 -88 -13887 88
rect -13763 -88 -13729 88
rect -13605 -88 -13571 88
rect -13447 -88 -13413 88
rect -13289 -88 -13255 88
rect -13131 -88 -13097 88
rect -12973 -88 -12939 88
rect -12815 -88 -12781 88
rect -12657 -88 -12623 88
rect -12499 -88 -12465 88
rect -12341 -88 -12307 88
rect -12183 -88 -12149 88
rect -12025 -88 -11991 88
rect -11867 -88 -11833 88
rect -11709 -88 -11675 88
rect -11551 -88 -11517 88
rect -11393 -88 -11359 88
rect -11235 -88 -11201 88
rect -11077 -88 -11043 88
rect -10919 -88 -10885 88
rect -10761 -88 -10727 88
rect -10603 -88 -10569 88
rect -10445 -88 -10411 88
rect -10287 -88 -10253 88
rect -10129 -88 -10095 88
rect -9971 -88 -9937 88
rect -9813 -88 -9779 88
rect -9655 -88 -9621 88
rect -9497 -88 -9463 88
rect -9339 -88 -9305 88
rect -9181 -88 -9147 88
rect -9023 -88 -8989 88
rect -8865 -88 -8831 88
rect -8707 -88 -8673 88
rect -8549 -88 -8515 88
rect -8391 -88 -8357 88
rect -8233 -88 -8199 88
rect -8075 -88 -8041 88
rect -7917 -88 -7883 88
rect -7759 -88 -7725 88
rect -7601 -88 -7567 88
rect -7443 -88 -7409 88
rect -7285 -88 -7251 88
rect -7127 -88 -7093 88
rect -6969 -88 -6935 88
rect -6811 -88 -6777 88
rect -6653 -88 -6619 88
rect -6495 -88 -6461 88
rect -6337 -88 -6303 88
rect -6179 -88 -6145 88
rect -6021 -88 -5987 88
rect -5863 -88 -5829 88
rect -5705 -88 -5671 88
rect -5547 -88 -5513 88
rect -5389 -88 -5355 88
rect -5231 -88 -5197 88
rect -5073 -88 -5039 88
rect -4915 -88 -4881 88
rect -4757 -88 -4723 88
rect -4599 -88 -4565 88
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect 4565 -88 4599 88
rect 4723 -88 4757 88
rect 4881 -88 4915 88
rect 5039 -88 5073 88
rect 5197 -88 5231 88
rect 5355 -88 5389 88
rect 5513 -88 5547 88
rect 5671 -88 5705 88
rect 5829 -88 5863 88
rect 5987 -88 6021 88
rect 6145 -88 6179 88
rect 6303 -88 6337 88
rect 6461 -88 6495 88
rect 6619 -88 6653 88
rect 6777 -88 6811 88
rect 6935 -88 6969 88
rect 7093 -88 7127 88
rect 7251 -88 7285 88
rect 7409 -88 7443 88
rect 7567 -88 7601 88
rect 7725 -88 7759 88
rect 7883 -88 7917 88
rect 8041 -88 8075 88
rect 8199 -88 8233 88
rect 8357 -88 8391 88
rect 8515 -88 8549 88
rect 8673 -88 8707 88
rect 8831 -88 8865 88
rect 8989 -88 9023 88
rect 9147 -88 9181 88
rect 9305 -88 9339 88
rect 9463 -88 9497 88
rect 9621 -88 9655 88
rect 9779 -88 9813 88
rect 9937 -88 9971 88
rect 10095 -88 10129 88
rect 10253 -88 10287 88
rect 10411 -88 10445 88
rect 10569 -88 10603 88
rect 10727 -88 10761 88
rect 10885 -88 10919 88
rect 11043 -88 11077 88
rect 11201 -88 11235 88
rect 11359 -88 11393 88
rect 11517 -88 11551 88
rect 11675 -88 11709 88
rect 11833 -88 11867 88
rect 11991 -88 12025 88
rect 12149 -88 12183 88
rect 12307 -88 12341 88
rect 12465 -88 12499 88
rect 12623 -88 12657 88
rect 12781 -88 12815 88
rect 12939 -88 12973 88
rect 13097 -88 13131 88
rect 13255 -88 13289 88
rect 13413 -88 13447 88
rect 13571 -88 13605 88
rect 13729 -88 13763 88
rect 13887 -88 13921 88
rect 14045 -88 14079 88
rect 14203 -88 14237 88
rect 14361 -88 14395 88
rect 14519 -88 14553 88
rect 14677 -88 14711 88
rect 14835 -88 14869 88
rect 14993 -88 15027 88
rect 15151 -88 15185 88
rect 15309 -88 15343 88
rect 15467 -88 15501 88
rect 15625 -88 15659 88
rect 15783 -88 15817 88
<< mvnsubdiff >>
rect -15963 319 15963 331
rect -15963 285 -15855 319
rect 15855 285 15963 319
rect -15963 273 15963 285
rect -15963 223 -15905 273
rect -15963 -223 -15951 223
rect -15917 -223 -15905 223
rect 15905 223 15963 273
rect -15963 -273 -15905 -223
rect 15905 -223 15917 223
rect 15951 -223 15963 223
rect 15905 -273 15963 -223
rect -15963 -285 15963 -273
rect -15963 -319 -15855 -285
rect 15855 -319 15963 -285
rect -15963 -331 15963 -319
<< mvnsubdiffcont >>
rect -15855 285 15855 319
rect -15951 -223 -15917 223
rect 15917 -223 15951 223
rect -15855 -319 15855 -285
<< poly >>
rect -15771 181 -15671 197
rect -15771 147 -15755 181
rect -15687 147 -15671 181
rect -15771 100 -15671 147
rect -15613 181 -15513 197
rect -15613 147 -15597 181
rect -15529 147 -15513 181
rect -15613 100 -15513 147
rect -15455 181 -15355 197
rect -15455 147 -15439 181
rect -15371 147 -15355 181
rect -15455 100 -15355 147
rect -15297 181 -15197 197
rect -15297 147 -15281 181
rect -15213 147 -15197 181
rect -15297 100 -15197 147
rect -15139 181 -15039 197
rect -15139 147 -15123 181
rect -15055 147 -15039 181
rect -15139 100 -15039 147
rect -14981 181 -14881 197
rect -14981 147 -14965 181
rect -14897 147 -14881 181
rect -14981 100 -14881 147
rect -14823 181 -14723 197
rect -14823 147 -14807 181
rect -14739 147 -14723 181
rect -14823 100 -14723 147
rect -14665 181 -14565 197
rect -14665 147 -14649 181
rect -14581 147 -14565 181
rect -14665 100 -14565 147
rect -14507 181 -14407 197
rect -14507 147 -14491 181
rect -14423 147 -14407 181
rect -14507 100 -14407 147
rect -14349 181 -14249 197
rect -14349 147 -14333 181
rect -14265 147 -14249 181
rect -14349 100 -14249 147
rect -14191 181 -14091 197
rect -14191 147 -14175 181
rect -14107 147 -14091 181
rect -14191 100 -14091 147
rect -14033 181 -13933 197
rect -14033 147 -14017 181
rect -13949 147 -13933 181
rect -14033 100 -13933 147
rect -13875 181 -13775 197
rect -13875 147 -13859 181
rect -13791 147 -13775 181
rect -13875 100 -13775 147
rect -13717 181 -13617 197
rect -13717 147 -13701 181
rect -13633 147 -13617 181
rect -13717 100 -13617 147
rect -13559 181 -13459 197
rect -13559 147 -13543 181
rect -13475 147 -13459 181
rect -13559 100 -13459 147
rect -13401 181 -13301 197
rect -13401 147 -13385 181
rect -13317 147 -13301 181
rect -13401 100 -13301 147
rect -13243 181 -13143 197
rect -13243 147 -13227 181
rect -13159 147 -13143 181
rect -13243 100 -13143 147
rect -13085 181 -12985 197
rect -13085 147 -13069 181
rect -13001 147 -12985 181
rect -13085 100 -12985 147
rect -12927 181 -12827 197
rect -12927 147 -12911 181
rect -12843 147 -12827 181
rect -12927 100 -12827 147
rect -12769 181 -12669 197
rect -12769 147 -12753 181
rect -12685 147 -12669 181
rect -12769 100 -12669 147
rect -12611 181 -12511 197
rect -12611 147 -12595 181
rect -12527 147 -12511 181
rect -12611 100 -12511 147
rect -12453 181 -12353 197
rect -12453 147 -12437 181
rect -12369 147 -12353 181
rect -12453 100 -12353 147
rect -12295 181 -12195 197
rect -12295 147 -12279 181
rect -12211 147 -12195 181
rect -12295 100 -12195 147
rect -12137 181 -12037 197
rect -12137 147 -12121 181
rect -12053 147 -12037 181
rect -12137 100 -12037 147
rect -11979 181 -11879 197
rect -11979 147 -11963 181
rect -11895 147 -11879 181
rect -11979 100 -11879 147
rect -11821 181 -11721 197
rect -11821 147 -11805 181
rect -11737 147 -11721 181
rect -11821 100 -11721 147
rect -11663 181 -11563 197
rect -11663 147 -11647 181
rect -11579 147 -11563 181
rect -11663 100 -11563 147
rect -11505 181 -11405 197
rect -11505 147 -11489 181
rect -11421 147 -11405 181
rect -11505 100 -11405 147
rect -11347 181 -11247 197
rect -11347 147 -11331 181
rect -11263 147 -11247 181
rect -11347 100 -11247 147
rect -11189 181 -11089 197
rect -11189 147 -11173 181
rect -11105 147 -11089 181
rect -11189 100 -11089 147
rect -11031 181 -10931 197
rect -11031 147 -11015 181
rect -10947 147 -10931 181
rect -11031 100 -10931 147
rect -10873 181 -10773 197
rect -10873 147 -10857 181
rect -10789 147 -10773 181
rect -10873 100 -10773 147
rect -10715 181 -10615 197
rect -10715 147 -10699 181
rect -10631 147 -10615 181
rect -10715 100 -10615 147
rect -10557 181 -10457 197
rect -10557 147 -10541 181
rect -10473 147 -10457 181
rect -10557 100 -10457 147
rect -10399 181 -10299 197
rect -10399 147 -10383 181
rect -10315 147 -10299 181
rect -10399 100 -10299 147
rect -10241 181 -10141 197
rect -10241 147 -10225 181
rect -10157 147 -10141 181
rect -10241 100 -10141 147
rect -10083 181 -9983 197
rect -10083 147 -10067 181
rect -9999 147 -9983 181
rect -10083 100 -9983 147
rect -9925 181 -9825 197
rect -9925 147 -9909 181
rect -9841 147 -9825 181
rect -9925 100 -9825 147
rect -9767 181 -9667 197
rect -9767 147 -9751 181
rect -9683 147 -9667 181
rect -9767 100 -9667 147
rect -9609 181 -9509 197
rect -9609 147 -9593 181
rect -9525 147 -9509 181
rect -9609 100 -9509 147
rect -9451 181 -9351 197
rect -9451 147 -9435 181
rect -9367 147 -9351 181
rect -9451 100 -9351 147
rect -9293 181 -9193 197
rect -9293 147 -9277 181
rect -9209 147 -9193 181
rect -9293 100 -9193 147
rect -9135 181 -9035 197
rect -9135 147 -9119 181
rect -9051 147 -9035 181
rect -9135 100 -9035 147
rect -8977 181 -8877 197
rect -8977 147 -8961 181
rect -8893 147 -8877 181
rect -8977 100 -8877 147
rect -8819 181 -8719 197
rect -8819 147 -8803 181
rect -8735 147 -8719 181
rect -8819 100 -8719 147
rect -8661 181 -8561 197
rect -8661 147 -8645 181
rect -8577 147 -8561 181
rect -8661 100 -8561 147
rect -8503 181 -8403 197
rect -8503 147 -8487 181
rect -8419 147 -8403 181
rect -8503 100 -8403 147
rect -8345 181 -8245 197
rect -8345 147 -8329 181
rect -8261 147 -8245 181
rect -8345 100 -8245 147
rect -8187 181 -8087 197
rect -8187 147 -8171 181
rect -8103 147 -8087 181
rect -8187 100 -8087 147
rect -8029 181 -7929 197
rect -8029 147 -8013 181
rect -7945 147 -7929 181
rect -8029 100 -7929 147
rect -7871 181 -7771 197
rect -7871 147 -7855 181
rect -7787 147 -7771 181
rect -7871 100 -7771 147
rect -7713 181 -7613 197
rect -7713 147 -7697 181
rect -7629 147 -7613 181
rect -7713 100 -7613 147
rect -7555 181 -7455 197
rect -7555 147 -7539 181
rect -7471 147 -7455 181
rect -7555 100 -7455 147
rect -7397 181 -7297 197
rect -7397 147 -7381 181
rect -7313 147 -7297 181
rect -7397 100 -7297 147
rect -7239 181 -7139 197
rect -7239 147 -7223 181
rect -7155 147 -7139 181
rect -7239 100 -7139 147
rect -7081 181 -6981 197
rect -7081 147 -7065 181
rect -6997 147 -6981 181
rect -7081 100 -6981 147
rect -6923 181 -6823 197
rect -6923 147 -6907 181
rect -6839 147 -6823 181
rect -6923 100 -6823 147
rect -6765 181 -6665 197
rect -6765 147 -6749 181
rect -6681 147 -6665 181
rect -6765 100 -6665 147
rect -6607 181 -6507 197
rect -6607 147 -6591 181
rect -6523 147 -6507 181
rect -6607 100 -6507 147
rect -6449 181 -6349 197
rect -6449 147 -6433 181
rect -6365 147 -6349 181
rect -6449 100 -6349 147
rect -6291 181 -6191 197
rect -6291 147 -6275 181
rect -6207 147 -6191 181
rect -6291 100 -6191 147
rect -6133 181 -6033 197
rect -6133 147 -6117 181
rect -6049 147 -6033 181
rect -6133 100 -6033 147
rect -5975 181 -5875 197
rect -5975 147 -5959 181
rect -5891 147 -5875 181
rect -5975 100 -5875 147
rect -5817 181 -5717 197
rect -5817 147 -5801 181
rect -5733 147 -5717 181
rect -5817 100 -5717 147
rect -5659 181 -5559 197
rect -5659 147 -5643 181
rect -5575 147 -5559 181
rect -5659 100 -5559 147
rect -5501 181 -5401 197
rect -5501 147 -5485 181
rect -5417 147 -5401 181
rect -5501 100 -5401 147
rect -5343 181 -5243 197
rect -5343 147 -5327 181
rect -5259 147 -5243 181
rect -5343 100 -5243 147
rect -5185 181 -5085 197
rect -5185 147 -5169 181
rect -5101 147 -5085 181
rect -5185 100 -5085 147
rect -5027 181 -4927 197
rect -5027 147 -5011 181
rect -4943 147 -4927 181
rect -5027 100 -4927 147
rect -4869 181 -4769 197
rect -4869 147 -4853 181
rect -4785 147 -4769 181
rect -4869 100 -4769 147
rect -4711 181 -4611 197
rect -4711 147 -4695 181
rect -4627 147 -4611 181
rect -4711 100 -4611 147
rect -4553 181 -4453 197
rect -4553 147 -4537 181
rect -4469 147 -4453 181
rect -4553 100 -4453 147
rect -4395 181 -4295 197
rect -4395 147 -4379 181
rect -4311 147 -4295 181
rect -4395 100 -4295 147
rect -4237 181 -4137 197
rect -4237 147 -4221 181
rect -4153 147 -4137 181
rect -4237 100 -4137 147
rect -4079 181 -3979 197
rect -4079 147 -4063 181
rect -3995 147 -3979 181
rect -4079 100 -3979 147
rect -3921 181 -3821 197
rect -3921 147 -3905 181
rect -3837 147 -3821 181
rect -3921 100 -3821 147
rect -3763 181 -3663 197
rect -3763 147 -3747 181
rect -3679 147 -3663 181
rect -3763 100 -3663 147
rect -3605 181 -3505 197
rect -3605 147 -3589 181
rect -3521 147 -3505 181
rect -3605 100 -3505 147
rect -3447 181 -3347 197
rect -3447 147 -3431 181
rect -3363 147 -3347 181
rect -3447 100 -3347 147
rect -3289 181 -3189 197
rect -3289 147 -3273 181
rect -3205 147 -3189 181
rect -3289 100 -3189 147
rect -3131 181 -3031 197
rect -3131 147 -3115 181
rect -3047 147 -3031 181
rect -3131 100 -3031 147
rect -2973 181 -2873 197
rect -2973 147 -2957 181
rect -2889 147 -2873 181
rect -2973 100 -2873 147
rect -2815 181 -2715 197
rect -2815 147 -2799 181
rect -2731 147 -2715 181
rect -2815 100 -2715 147
rect -2657 181 -2557 197
rect -2657 147 -2641 181
rect -2573 147 -2557 181
rect -2657 100 -2557 147
rect -2499 181 -2399 197
rect -2499 147 -2483 181
rect -2415 147 -2399 181
rect -2499 100 -2399 147
rect -2341 181 -2241 197
rect -2341 147 -2325 181
rect -2257 147 -2241 181
rect -2341 100 -2241 147
rect -2183 181 -2083 197
rect -2183 147 -2167 181
rect -2099 147 -2083 181
rect -2183 100 -2083 147
rect -2025 181 -1925 197
rect -2025 147 -2009 181
rect -1941 147 -1925 181
rect -2025 100 -1925 147
rect -1867 181 -1767 197
rect -1867 147 -1851 181
rect -1783 147 -1767 181
rect -1867 100 -1767 147
rect -1709 181 -1609 197
rect -1709 147 -1693 181
rect -1625 147 -1609 181
rect -1709 100 -1609 147
rect -1551 181 -1451 197
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1551 100 -1451 147
rect -1393 181 -1293 197
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1393 100 -1293 147
rect -1235 181 -1135 197
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1235 100 -1135 147
rect -1077 181 -977 197
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -1077 100 -977 147
rect -919 181 -819 197
rect -919 147 -903 181
rect -835 147 -819 181
rect -919 100 -819 147
rect -761 181 -661 197
rect -761 147 -745 181
rect -677 147 -661 181
rect -761 100 -661 147
rect -603 181 -503 197
rect -603 147 -587 181
rect -519 147 -503 181
rect -603 100 -503 147
rect -445 181 -345 197
rect -445 147 -429 181
rect -361 147 -345 181
rect -445 100 -345 147
rect -287 181 -187 197
rect -287 147 -271 181
rect -203 147 -187 181
rect -287 100 -187 147
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect 187 181 287 197
rect 187 147 203 181
rect 271 147 287 181
rect 187 100 287 147
rect 345 181 445 197
rect 345 147 361 181
rect 429 147 445 181
rect 345 100 445 147
rect 503 181 603 197
rect 503 147 519 181
rect 587 147 603 181
rect 503 100 603 147
rect 661 181 761 197
rect 661 147 677 181
rect 745 147 761 181
rect 661 100 761 147
rect 819 181 919 197
rect 819 147 835 181
rect 903 147 919 181
rect 819 100 919 147
rect 977 181 1077 197
rect 977 147 993 181
rect 1061 147 1077 181
rect 977 100 1077 147
rect 1135 181 1235 197
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1135 100 1235 147
rect 1293 181 1393 197
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1293 100 1393 147
rect 1451 181 1551 197
rect 1451 147 1467 181
rect 1535 147 1551 181
rect 1451 100 1551 147
rect 1609 181 1709 197
rect 1609 147 1625 181
rect 1693 147 1709 181
rect 1609 100 1709 147
rect 1767 181 1867 197
rect 1767 147 1783 181
rect 1851 147 1867 181
rect 1767 100 1867 147
rect 1925 181 2025 197
rect 1925 147 1941 181
rect 2009 147 2025 181
rect 1925 100 2025 147
rect 2083 181 2183 197
rect 2083 147 2099 181
rect 2167 147 2183 181
rect 2083 100 2183 147
rect 2241 181 2341 197
rect 2241 147 2257 181
rect 2325 147 2341 181
rect 2241 100 2341 147
rect 2399 181 2499 197
rect 2399 147 2415 181
rect 2483 147 2499 181
rect 2399 100 2499 147
rect 2557 181 2657 197
rect 2557 147 2573 181
rect 2641 147 2657 181
rect 2557 100 2657 147
rect 2715 181 2815 197
rect 2715 147 2731 181
rect 2799 147 2815 181
rect 2715 100 2815 147
rect 2873 181 2973 197
rect 2873 147 2889 181
rect 2957 147 2973 181
rect 2873 100 2973 147
rect 3031 181 3131 197
rect 3031 147 3047 181
rect 3115 147 3131 181
rect 3031 100 3131 147
rect 3189 181 3289 197
rect 3189 147 3205 181
rect 3273 147 3289 181
rect 3189 100 3289 147
rect 3347 181 3447 197
rect 3347 147 3363 181
rect 3431 147 3447 181
rect 3347 100 3447 147
rect 3505 181 3605 197
rect 3505 147 3521 181
rect 3589 147 3605 181
rect 3505 100 3605 147
rect 3663 181 3763 197
rect 3663 147 3679 181
rect 3747 147 3763 181
rect 3663 100 3763 147
rect 3821 181 3921 197
rect 3821 147 3837 181
rect 3905 147 3921 181
rect 3821 100 3921 147
rect 3979 181 4079 197
rect 3979 147 3995 181
rect 4063 147 4079 181
rect 3979 100 4079 147
rect 4137 181 4237 197
rect 4137 147 4153 181
rect 4221 147 4237 181
rect 4137 100 4237 147
rect 4295 181 4395 197
rect 4295 147 4311 181
rect 4379 147 4395 181
rect 4295 100 4395 147
rect 4453 181 4553 197
rect 4453 147 4469 181
rect 4537 147 4553 181
rect 4453 100 4553 147
rect 4611 181 4711 197
rect 4611 147 4627 181
rect 4695 147 4711 181
rect 4611 100 4711 147
rect 4769 181 4869 197
rect 4769 147 4785 181
rect 4853 147 4869 181
rect 4769 100 4869 147
rect 4927 181 5027 197
rect 4927 147 4943 181
rect 5011 147 5027 181
rect 4927 100 5027 147
rect 5085 181 5185 197
rect 5085 147 5101 181
rect 5169 147 5185 181
rect 5085 100 5185 147
rect 5243 181 5343 197
rect 5243 147 5259 181
rect 5327 147 5343 181
rect 5243 100 5343 147
rect 5401 181 5501 197
rect 5401 147 5417 181
rect 5485 147 5501 181
rect 5401 100 5501 147
rect 5559 181 5659 197
rect 5559 147 5575 181
rect 5643 147 5659 181
rect 5559 100 5659 147
rect 5717 181 5817 197
rect 5717 147 5733 181
rect 5801 147 5817 181
rect 5717 100 5817 147
rect 5875 181 5975 197
rect 5875 147 5891 181
rect 5959 147 5975 181
rect 5875 100 5975 147
rect 6033 181 6133 197
rect 6033 147 6049 181
rect 6117 147 6133 181
rect 6033 100 6133 147
rect 6191 181 6291 197
rect 6191 147 6207 181
rect 6275 147 6291 181
rect 6191 100 6291 147
rect 6349 181 6449 197
rect 6349 147 6365 181
rect 6433 147 6449 181
rect 6349 100 6449 147
rect 6507 181 6607 197
rect 6507 147 6523 181
rect 6591 147 6607 181
rect 6507 100 6607 147
rect 6665 181 6765 197
rect 6665 147 6681 181
rect 6749 147 6765 181
rect 6665 100 6765 147
rect 6823 181 6923 197
rect 6823 147 6839 181
rect 6907 147 6923 181
rect 6823 100 6923 147
rect 6981 181 7081 197
rect 6981 147 6997 181
rect 7065 147 7081 181
rect 6981 100 7081 147
rect 7139 181 7239 197
rect 7139 147 7155 181
rect 7223 147 7239 181
rect 7139 100 7239 147
rect 7297 181 7397 197
rect 7297 147 7313 181
rect 7381 147 7397 181
rect 7297 100 7397 147
rect 7455 181 7555 197
rect 7455 147 7471 181
rect 7539 147 7555 181
rect 7455 100 7555 147
rect 7613 181 7713 197
rect 7613 147 7629 181
rect 7697 147 7713 181
rect 7613 100 7713 147
rect 7771 181 7871 197
rect 7771 147 7787 181
rect 7855 147 7871 181
rect 7771 100 7871 147
rect 7929 181 8029 197
rect 7929 147 7945 181
rect 8013 147 8029 181
rect 7929 100 8029 147
rect 8087 181 8187 197
rect 8087 147 8103 181
rect 8171 147 8187 181
rect 8087 100 8187 147
rect 8245 181 8345 197
rect 8245 147 8261 181
rect 8329 147 8345 181
rect 8245 100 8345 147
rect 8403 181 8503 197
rect 8403 147 8419 181
rect 8487 147 8503 181
rect 8403 100 8503 147
rect 8561 181 8661 197
rect 8561 147 8577 181
rect 8645 147 8661 181
rect 8561 100 8661 147
rect 8719 181 8819 197
rect 8719 147 8735 181
rect 8803 147 8819 181
rect 8719 100 8819 147
rect 8877 181 8977 197
rect 8877 147 8893 181
rect 8961 147 8977 181
rect 8877 100 8977 147
rect 9035 181 9135 197
rect 9035 147 9051 181
rect 9119 147 9135 181
rect 9035 100 9135 147
rect 9193 181 9293 197
rect 9193 147 9209 181
rect 9277 147 9293 181
rect 9193 100 9293 147
rect 9351 181 9451 197
rect 9351 147 9367 181
rect 9435 147 9451 181
rect 9351 100 9451 147
rect 9509 181 9609 197
rect 9509 147 9525 181
rect 9593 147 9609 181
rect 9509 100 9609 147
rect 9667 181 9767 197
rect 9667 147 9683 181
rect 9751 147 9767 181
rect 9667 100 9767 147
rect 9825 181 9925 197
rect 9825 147 9841 181
rect 9909 147 9925 181
rect 9825 100 9925 147
rect 9983 181 10083 197
rect 9983 147 9999 181
rect 10067 147 10083 181
rect 9983 100 10083 147
rect 10141 181 10241 197
rect 10141 147 10157 181
rect 10225 147 10241 181
rect 10141 100 10241 147
rect 10299 181 10399 197
rect 10299 147 10315 181
rect 10383 147 10399 181
rect 10299 100 10399 147
rect 10457 181 10557 197
rect 10457 147 10473 181
rect 10541 147 10557 181
rect 10457 100 10557 147
rect 10615 181 10715 197
rect 10615 147 10631 181
rect 10699 147 10715 181
rect 10615 100 10715 147
rect 10773 181 10873 197
rect 10773 147 10789 181
rect 10857 147 10873 181
rect 10773 100 10873 147
rect 10931 181 11031 197
rect 10931 147 10947 181
rect 11015 147 11031 181
rect 10931 100 11031 147
rect 11089 181 11189 197
rect 11089 147 11105 181
rect 11173 147 11189 181
rect 11089 100 11189 147
rect 11247 181 11347 197
rect 11247 147 11263 181
rect 11331 147 11347 181
rect 11247 100 11347 147
rect 11405 181 11505 197
rect 11405 147 11421 181
rect 11489 147 11505 181
rect 11405 100 11505 147
rect 11563 181 11663 197
rect 11563 147 11579 181
rect 11647 147 11663 181
rect 11563 100 11663 147
rect 11721 181 11821 197
rect 11721 147 11737 181
rect 11805 147 11821 181
rect 11721 100 11821 147
rect 11879 181 11979 197
rect 11879 147 11895 181
rect 11963 147 11979 181
rect 11879 100 11979 147
rect 12037 181 12137 197
rect 12037 147 12053 181
rect 12121 147 12137 181
rect 12037 100 12137 147
rect 12195 181 12295 197
rect 12195 147 12211 181
rect 12279 147 12295 181
rect 12195 100 12295 147
rect 12353 181 12453 197
rect 12353 147 12369 181
rect 12437 147 12453 181
rect 12353 100 12453 147
rect 12511 181 12611 197
rect 12511 147 12527 181
rect 12595 147 12611 181
rect 12511 100 12611 147
rect 12669 181 12769 197
rect 12669 147 12685 181
rect 12753 147 12769 181
rect 12669 100 12769 147
rect 12827 181 12927 197
rect 12827 147 12843 181
rect 12911 147 12927 181
rect 12827 100 12927 147
rect 12985 181 13085 197
rect 12985 147 13001 181
rect 13069 147 13085 181
rect 12985 100 13085 147
rect 13143 181 13243 197
rect 13143 147 13159 181
rect 13227 147 13243 181
rect 13143 100 13243 147
rect 13301 181 13401 197
rect 13301 147 13317 181
rect 13385 147 13401 181
rect 13301 100 13401 147
rect 13459 181 13559 197
rect 13459 147 13475 181
rect 13543 147 13559 181
rect 13459 100 13559 147
rect 13617 181 13717 197
rect 13617 147 13633 181
rect 13701 147 13717 181
rect 13617 100 13717 147
rect 13775 181 13875 197
rect 13775 147 13791 181
rect 13859 147 13875 181
rect 13775 100 13875 147
rect 13933 181 14033 197
rect 13933 147 13949 181
rect 14017 147 14033 181
rect 13933 100 14033 147
rect 14091 181 14191 197
rect 14091 147 14107 181
rect 14175 147 14191 181
rect 14091 100 14191 147
rect 14249 181 14349 197
rect 14249 147 14265 181
rect 14333 147 14349 181
rect 14249 100 14349 147
rect 14407 181 14507 197
rect 14407 147 14423 181
rect 14491 147 14507 181
rect 14407 100 14507 147
rect 14565 181 14665 197
rect 14565 147 14581 181
rect 14649 147 14665 181
rect 14565 100 14665 147
rect 14723 181 14823 197
rect 14723 147 14739 181
rect 14807 147 14823 181
rect 14723 100 14823 147
rect 14881 181 14981 197
rect 14881 147 14897 181
rect 14965 147 14981 181
rect 14881 100 14981 147
rect 15039 181 15139 197
rect 15039 147 15055 181
rect 15123 147 15139 181
rect 15039 100 15139 147
rect 15197 181 15297 197
rect 15197 147 15213 181
rect 15281 147 15297 181
rect 15197 100 15297 147
rect 15355 181 15455 197
rect 15355 147 15371 181
rect 15439 147 15455 181
rect 15355 100 15455 147
rect 15513 181 15613 197
rect 15513 147 15529 181
rect 15597 147 15613 181
rect 15513 100 15613 147
rect 15671 181 15771 197
rect 15671 147 15687 181
rect 15755 147 15771 181
rect 15671 100 15771 147
rect -15771 -147 -15671 -100
rect -15771 -181 -15755 -147
rect -15687 -181 -15671 -147
rect -15771 -197 -15671 -181
rect -15613 -147 -15513 -100
rect -15613 -181 -15597 -147
rect -15529 -181 -15513 -147
rect -15613 -197 -15513 -181
rect -15455 -147 -15355 -100
rect -15455 -181 -15439 -147
rect -15371 -181 -15355 -147
rect -15455 -197 -15355 -181
rect -15297 -147 -15197 -100
rect -15297 -181 -15281 -147
rect -15213 -181 -15197 -147
rect -15297 -197 -15197 -181
rect -15139 -147 -15039 -100
rect -15139 -181 -15123 -147
rect -15055 -181 -15039 -147
rect -15139 -197 -15039 -181
rect -14981 -147 -14881 -100
rect -14981 -181 -14965 -147
rect -14897 -181 -14881 -147
rect -14981 -197 -14881 -181
rect -14823 -147 -14723 -100
rect -14823 -181 -14807 -147
rect -14739 -181 -14723 -147
rect -14823 -197 -14723 -181
rect -14665 -147 -14565 -100
rect -14665 -181 -14649 -147
rect -14581 -181 -14565 -147
rect -14665 -197 -14565 -181
rect -14507 -147 -14407 -100
rect -14507 -181 -14491 -147
rect -14423 -181 -14407 -147
rect -14507 -197 -14407 -181
rect -14349 -147 -14249 -100
rect -14349 -181 -14333 -147
rect -14265 -181 -14249 -147
rect -14349 -197 -14249 -181
rect -14191 -147 -14091 -100
rect -14191 -181 -14175 -147
rect -14107 -181 -14091 -147
rect -14191 -197 -14091 -181
rect -14033 -147 -13933 -100
rect -14033 -181 -14017 -147
rect -13949 -181 -13933 -147
rect -14033 -197 -13933 -181
rect -13875 -147 -13775 -100
rect -13875 -181 -13859 -147
rect -13791 -181 -13775 -147
rect -13875 -197 -13775 -181
rect -13717 -147 -13617 -100
rect -13717 -181 -13701 -147
rect -13633 -181 -13617 -147
rect -13717 -197 -13617 -181
rect -13559 -147 -13459 -100
rect -13559 -181 -13543 -147
rect -13475 -181 -13459 -147
rect -13559 -197 -13459 -181
rect -13401 -147 -13301 -100
rect -13401 -181 -13385 -147
rect -13317 -181 -13301 -147
rect -13401 -197 -13301 -181
rect -13243 -147 -13143 -100
rect -13243 -181 -13227 -147
rect -13159 -181 -13143 -147
rect -13243 -197 -13143 -181
rect -13085 -147 -12985 -100
rect -13085 -181 -13069 -147
rect -13001 -181 -12985 -147
rect -13085 -197 -12985 -181
rect -12927 -147 -12827 -100
rect -12927 -181 -12911 -147
rect -12843 -181 -12827 -147
rect -12927 -197 -12827 -181
rect -12769 -147 -12669 -100
rect -12769 -181 -12753 -147
rect -12685 -181 -12669 -147
rect -12769 -197 -12669 -181
rect -12611 -147 -12511 -100
rect -12611 -181 -12595 -147
rect -12527 -181 -12511 -147
rect -12611 -197 -12511 -181
rect -12453 -147 -12353 -100
rect -12453 -181 -12437 -147
rect -12369 -181 -12353 -147
rect -12453 -197 -12353 -181
rect -12295 -147 -12195 -100
rect -12295 -181 -12279 -147
rect -12211 -181 -12195 -147
rect -12295 -197 -12195 -181
rect -12137 -147 -12037 -100
rect -12137 -181 -12121 -147
rect -12053 -181 -12037 -147
rect -12137 -197 -12037 -181
rect -11979 -147 -11879 -100
rect -11979 -181 -11963 -147
rect -11895 -181 -11879 -147
rect -11979 -197 -11879 -181
rect -11821 -147 -11721 -100
rect -11821 -181 -11805 -147
rect -11737 -181 -11721 -147
rect -11821 -197 -11721 -181
rect -11663 -147 -11563 -100
rect -11663 -181 -11647 -147
rect -11579 -181 -11563 -147
rect -11663 -197 -11563 -181
rect -11505 -147 -11405 -100
rect -11505 -181 -11489 -147
rect -11421 -181 -11405 -147
rect -11505 -197 -11405 -181
rect -11347 -147 -11247 -100
rect -11347 -181 -11331 -147
rect -11263 -181 -11247 -147
rect -11347 -197 -11247 -181
rect -11189 -147 -11089 -100
rect -11189 -181 -11173 -147
rect -11105 -181 -11089 -147
rect -11189 -197 -11089 -181
rect -11031 -147 -10931 -100
rect -11031 -181 -11015 -147
rect -10947 -181 -10931 -147
rect -11031 -197 -10931 -181
rect -10873 -147 -10773 -100
rect -10873 -181 -10857 -147
rect -10789 -181 -10773 -147
rect -10873 -197 -10773 -181
rect -10715 -147 -10615 -100
rect -10715 -181 -10699 -147
rect -10631 -181 -10615 -147
rect -10715 -197 -10615 -181
rect -10557 -147 -10457 -100
rect -10557 -181 -10541 -147
rect -10473 -181 -10457 -147
rect -10557 -197 -10457 -181
rect -10399 -147 -10299 -100
rect -10399 -181 -10383 -147
rect -10315 -181 -10299 -147
rect -10399 -197 -10299 -181
rect -10241 -147 -10141 -100
rect -10241 -181 -10225 -147
rect -10157 -181 -10141 -147
rect -10241 -197 -10141 -181
rect -10083 -147 -9983 -100
rect -10083 -181 -10067 -147
rect -9999 -181 -9983 -147
rect -10083 -197 -9983 -181
rect -9925 -147 -9825 -100
rect -9925 -181 -9909 -147
rect -9841 -181 -9825 -147
rect -9925 -197 -9825 -181
rect -9767 -147 -9667 -100
rect -9767 -181 -9751 -147
rect -9683 -181 -9667 -147
rect -9767 -197 -9667 -181
rect -9609 -147 -9509 -100
rect -9609 -181 -9593 -147
rect -9525 -181 -9509 -147
rect -9609 -197 -9509 -181
rect -9451 -147 -9351 -100
rect -9451 -181 -9435 -147
rect -9367 -181 -9351 -147
rect -9451 -197 -9351 -181
rect -9293 -147 -9193 -100
rect -9293 -181 -9277 -147
rect -9209 -181 -9193 -147
rect -9293 -197 -9193 -181
rect -9135 -147 -9035 -100
rect -9135 -181 -9119 -147
rect -9051 -181 -9035 -147
rect -9135 -197 -9035 -181
rect -8977 -147 -8877 -100
rect -8977 -181 -8961 -147
rect -8893 -181 -8877 -147
rect -8977 -197 -8877 -181
rect -8819 -147 -8719 -100
rect -8819 -181 -8803 -147
rect -8735 -181 -8719 -147
rect -8819 -197 -8719 -181
rect -8661 -147 -8561 -100
rect -8661 -181 -8645 -147
rect -8577 -181 -8561 -147
rect -8661 -197 -8561 -181
rect -8503 -147 -8403 -100
rect -8503 -181 -8487 -147
rect -8419 -181 -8403 -147
rect -8503 -197 -8403 -181
rect -8345 -147 -8245 -100
rect -8345 -181 -8329 -147
rect -8261 -181 -8245 -147
rect -8345 -197 -8245 -181
rect -8187 -147 -8087 -100
rect -8187 -181 -8171 -147
rect -8103 -181 -8087 -147
rect -8187 -197 -8087 -181
rect -8029 -147 -7929 -100
rect -8029 -181 -8013 -147
rect -7945 -181 -7929 -147
rect -8029 -197 -7929 -181
rect -7871 -147 -7771 -100
rect -7871 -181 -7855 -147
rect -7787 -181 -7771 -147
rect -7871 -197 -7771 -181
rect -7713 -147 -7613 -100
rect -7713 -181 -7697 -147
rect -7629 -181 -7613 -147
rect -7713 -197 -7613 -181
rect -7555 -147 -7455 -100
rect -7555 -181 -7539 -147
rect -7471 -181 -7455 -147
rect -7555 -197 -7455 -181
rect -7397 -147 -7297 -100
rect -7397 -181 -7381 -147
rect -7313 -181 -7297 -147
rect -7397 -197 -7297 -181
rect -7239 -147 -7139 -100
rect -7239 -181 -7223 -147
rect -7155 -181 -7139 -147
rect -7239 -197 -7139 -181
rect -7081 -147 -6981 -100
rect -7081 -181 -7065 -147
rect -6997 -181 -6981 -147
rect -7081 -197 -6981 -181
rect -6923 -147 -6823 -100
rect -6923 -181 -6907 -147
rect -6839 -181 -6823 -147
rect -6923 -197 -6823 -181
rect -6765 -147 -6665 -100
rect -6765 -181 -6749 -147
rect -6681 -181 -6665 -147
rect -6765 -197 -6665 -181
rect -6607 -147 -6507 -100
rect -6607 -181 -6591 -147
rect -6523 -181 -6507 -147
rect -6607 -197 -6507 -181
rect -6449 -147 -6349 -100
rect -6449 -181 -6433 -147
rect -6365 -181 -6349 -147
rect -6449 -197 -6349 -181
rect -6291 -147 -6191 -100
rect -6291 -181 -6275 -147
rect -6207 -181 -6191 -147
rect -6291 -197 -6191 -181
rect -6133 -147 -6033 -100
rect -6133 -181 -6117 -147
rect -6049 -181 -6033 -147
rect -6133 -197 -6033 -181
rect -5975 -147 -5875 -100
rect -5975 -181 -5959 -147
rect -5891 -181 -5875 -147
rect -5975 -197 -5875 -181
rect -5817 -147 -5717 -100
rect -5817 -181 -5801 -147
rect -5733 -181 -5717 -147
rect -5817 -197 -5717 -181
rect -5659 -147 -5559 -100
rect -5659 -181 -5643 -147
rect -5575 -181 -5559 -147
rect -5659 -197 -5559 -181
rect -5501 -147 -5401 -100
rect -5501 -181 -5485 -147
rect -5417 -181 -5401 -147
rect -5501 -197 -5401 -181
rect -5343 -147 -5243 -100
rect -5343 -181 -5327 -147
rect -5259 -181 -5243 -147
rect -5343 -197 -5243 -181
rect -5185 -147 -5085 -100
rect -5185 -181 -5169 -147
rect -5101 -181 -5085 -147
rect -5185 -197 -5085 -181
rect -5027 -147 -4927 -100
rect -5027 -181 -5011 -147
rect -4943 -181 -4927 -147
rect -5027 -197 -4927 -181
rect -4869 -147 -4769 -100
rect -4869 -181 -4853 -147
rect -4785 -181 -4769 -147
rect -4869 -197 -4769 -181
rect -4711 -147 -4611 -100
rect -4711 -181 -4695 -147
rect -4627 -181 -4611 -147
rect -4711 -197 -4611 -181
rect -4553 -147 -4453 -100
rect -4553 -181 -4537 -147
rect -4469 -181 -4453 -147
rect -4553 -197 -4453 -181
rect -4395 -147 -4295 -100
rect -4395 -181 -4379 -147
rect -4311 -181 -4295 -147
rect -4395 -197 -4295 -181
rect -4237 -147 -4137 -100
rect -4237 -181 -4221 -147
rect -4153 -181 -4137 -147
rect -4237 -197 -4137 -181
rect -4079 -147 -3979 -100
rect -4079 -181 -4063 -147
rect -3995 -181 -3979 -147
rect -4079 -197 -3979 -181
rect -3921 -147 -3821 -100
rect -3921 -181 -3905 -147
rect -3837 -181 -3821 -147
rect -3921 -197 -3821 -181
rect -3763 -147 -3663 -100
rect -3763 -181 -3747 -147
rect -3679 -181 -3663 -147
rect -3763 -197 -3663 -181
rect -3605 -147 -3505 -100
rect -3605 -181 -3589 -147
rect -3521 -181 -3505 -147
rect -3605 -197 -3505 -181
rect -3447 -147 -3347 -100
rect -3447 -181 -3431 -147
rect -3363 -181 -3347 -147
rect -3447 -197 -3347 -181
rect -3289 -147 -3189 -100
rect -3289 -181 -3273 -147
rect -3205 -181 -3189 -147
rect -3289 -197 -3189 -181
rect -3131 -147 -3031 -100
rect -3131 -181 -3115 -147
rect -3047 -181 -3031 -147
rect -3131 -197 -3031 -181
rect -2973 -147 -2873 -100
rect -2973 -181 -2957 -147
rect -2889 -181 -2873 -147
rect -2973 -197 -2873 -181
rect -2815 -147 -2715 -100
rect -2815 -181 -2799 -147
rect -2731 -181 -2715 -147
rect -2815 -197 -2715 -181
rect -2657 -147 -2557 -100
rect -2657 -181 -2641 -147
rect -2573 -181 -2557 -147
rect -2657 -197 -2557 -181
rect -2499 -147 -2399 -100
rect -2499 -181 -2483 -147
rect -2415 -181 -2399 -147
rect -2499 -197 -2399 -181
rect -2341 -147 -2241 -100
rect -2341 -181 -2325 -147
rect -2257 -181 -2241 -147
rect -2341 -197 -2241 -181
rect -2183 -147 -2083 -100
rect -2183 -181 -2167 -147
rect -2099 -181 -2083 -147
rect -2183 -197 -2083 -181
rect -2025 -147 -1925 -100
rect -2025 -181 -2009 -147
rect -1941 -181 -1925 -147
rect -2025 -197 -1925 -181
rect -1867 -147 -1767 -100
rect -1867 -181 -1851 -147
rect -1783 -181 -1767 -147
rect -1867 -197 -1767 -181
rect -1709 -147 -1609 -100
rect -1709 -181 -1693 -147
rect -1625 -181 -1609 -147
rect -1709 -197 -1609 -181
rect -1551 -147 -1451 -100
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1551 -197 -1451 -181
rect -1393 -147 -1293 -100
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1393 -197 -1293 -181
rect -1235 -147 -1135 -100
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1235 -197 -1135 -181
rect -1077 -147 -977 -100
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -1077 -197 -977 -181
rect -919 -147 -819 -100
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -919 -197 -819 -181
rect -761 -147 -661 -100
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -761 -197 -661 -181
rect -603 -147 -503 -100
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -603 -197 -503 -181
rect -445 -147 -345 -100
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -445 -197 -345 -181
rect -287 -147 -187 -100
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -287 -197 -187 -181
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
rect 187 -147 287 -100
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 187 -197 287 -181
rect 345 -147 445 -100
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 345 -197 445 -181
rect 503 -147 603 -100
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 503 -197 603 -181
rect 661 -147 761 -100
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 661 -197 761 -181
rect 819 -147 919 -100
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 819 -197 919 -181
rect 977 -147 1077 -100
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 977 -197 1077 -181
rect 1135 -147 1235 -100
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1135 -197 1235 -181
rect 1293 -147 1393 -100
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1293 -197 1393 -181
rect 1451 -147 1551 -100
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect 1451 -197 1551 -181
rect 1609 -147 1709 -100
rect 1609 -181 1625 -147
rect 1693 -181 1709 -147
rect 1609 -197 1709 -181
rect 1767 -147 1867 -100
rect 1767 -181 1783 -147
rect 1851 -181 1867 -147
rect 1767 -197 1867 -181
rect 1925 -147 2025 -100
rect 1925 -181 1941 -147
rect 2009 -181 2025 -147
rect 1925 -197 2025 -181
rect 2083 -147 2183 -100
rect 2083 -181 2099 -147
rect 2167 -181 2183 -147
rect 2083 -197 2183 -181
rect 2241 -147 2341 -100
rect 2241 -181 2257 -147
rect 2325 -181 2341 -147
rect 2241 -197 2341 -181
rect 2399 -147 2499 -100
rect 2399 -181 2415 -147
rect 2483 -181 2499 -147
rect 2399 -197 2499 -181
rect 2557 -147 2657 -100
rect 2557 -181 2573 -147
rect 2641 -181 2657 -147
rect 2557 -197 2657 -181
rect 2715 -147 2815 -100
rect 2715 -181 2731 -147
rect 2799 -181 2815 -147
rect 2715 -197 2815 -181
rect 2873 -147 2973 -100
rect 2873 -181 2889 -147
rect 2957 -181 2973 -147
rect 2873 -197 2973 -181
rect 3031 -147 3131 -100
rect 3031 -181 3047 -147
rect 3115 -181 3131 -147
rect 3031 -197 3131 -181
rect 3189 -147 3289 -100
rect 3189 -181 3205 -147
rect 3273 -181 3289 -147
rect 3189 -197 3289 -181
rect 3347 -147 3447 -100
rect 3347 -181 3363 -147
rect 3431 -181 3447 -147
rect 3347 -197 3447 -181
rect 3505 -147 3605 -100
rect 3505 -181 3521 -147
rect 3589 -181 3605 -147
rect 3505 -197 3605 -181
rect 3663 -147 3763 -100
rect 3663 -181 3679 -147
rect 3747 -181 3763 -147
rect 3663 -197 3763 -181
rect 3821 -147 3921 -100
rect 3821 -181 3837 -147
rect 3905 -181 3921 -147
rect 3821 -197 3921 -181
rect 3979 -147 4079 -100
rect 3979 -181 3995 -147
rect 4063 -181 4079 -147
rect 3979 -197 4079 -181
rect 4137 -147 4237 -100
rect 4137 -181 4153 -147
rect 4221 -181 4237 -147
rect 4137 -197 4237 -181
rect 4295 -147 4395 -100
rect 4295 -181 4311 -147
rect 4379 -181 4395 -147
rect 4295 -197 4395 -181
rect 4453 -147 4553 -100
rect 4453 -181 4469 -147
rect 4537 -181 4553 -147
rect 4453 -197 4553 -181
rect 4611 -147 4711 -100
rect 4611 -181 4627 -147
rect 4695 -181 4711 -147
rect 4611 -197 4711 -181
rect 4769 -147 4869 -100
rect 4769 -181 4785 -147
rect 4853 -181 4869 -147
rect 4769 -197 4869 -181
rect 4927 -147 5027 -100
rect 4927 -181 4943 -147
rect 5011 -181 5027 -147
rect 4927 -197 5027 -181
rect 5085 -147 5185 -100
rect 5085 -181 5101 -147
rect 5169 -181 5185 -147
rect 5085 -197 5185 -181
rect 5243 -147 5343 -100
rect 5243 -181 5259 -147
rect 5327 -181 5343 -147
rect 5243 -197 5343 -181
rect 5401 -147 5501 -100
rect 5401 -181 5417 -147
rect 5485 -181 5501 -147
rect 5401 -197 5501 -181
rect 5559 -147 5659 -100
rect 5559 -181 5575 -147
rect 5643 -181 5659 -147
rect 5559 -197 5659 -181
rect 5717 -147 5817 -100
rect 5717 -181 5733 -147
rect 5801 -181 5817 -147
rect 5717 -197 5817 -181
rect 5875 -147 5975 -100
rect 5875 -181 5891 -147
rect 5959 -181 5975 -147
rect 5875 -197 5975 -181
rect 6033 -147 6133 -100
rect 6033 -181 6049 -147
rect 6117 -181 6133 -147
rect 6033 -197 6133 -181
rect 6191 -147 6291 -100
rect 6191 -181 6207 -147
rect 6275 -181 6291 -147
rect 6191 -197 6291 -181
rect 6349 -147 6449 -100
rect 6349 -181 6365 -147
rect 6433 -181 6449 -147
rect 6349 -197 6449 -181
rect 6507 -147 6607 -100
rect 6507 -181 6523 -147
rect 6591 -181 6607 -147
rect 6507 -197 6607 -181
rect 6665 -147 6765 -100
rect 6665 -181 6681 -147
rect 6749 -181 6765 -147
rect 6665 -197 6765 -181
rect 6823 -147 6923 -100
rect 6823 -181 6839 -147
rect 6907 -181 6923 -147
rect 6823 -197 6923 -181
rect 6981 -147 7081 -100
rect 6981 -181 6997 -147
rect 7065 -181 7081 -147
rect 6981 -197 7081 -181
rect 7139 -147 7239 -100
rect 7139 -181 7155 -147
rect 7223 -181 7239 -147
rect 7139 -197 7239 -181
rect 7297 -147 7397 -100
rect 7297 -181 7313 -147
rect 7381 -181 7397 -147
rect 7297 -197 7397 -181
rect 7455 -147 7555 -100
rect 7455 -181 7471 -147
rect 7539 -181 7555 -147
rect 7455 -197 7555 -181
rect 7613 -147 7713 -100
rect 7613 -181 7629 -147
rect 7697 -181 7713 -147
rect 7613 -197 7713 -181
rect 7771 -147 7871 -100
rect 7771 -181 7787 -147
rect 7855 -181 7871 -147
rect 7771 -197 7871 -181
rect 7929 -147 8029 -100
rect 7929 -181 7945 -147
rect 8013 -181 8029 -147
rect 7929 -197 8029 -181
rect 8087 -147 8187 -100
rect 8087 -181 8103 -147
rect 8171 -181 8187 -147
rect 8087 -197 8187 -181
rect 8245 -147 8345 -100
rect 8245 -181 8261 -147
rect 8329 -181 8345 -147
rect 8245 -197 8345 -181
rect 8403 -147 8503 -100
rect 8403 -181 8419 -147
rect 8487 -181 8503 -147
rect 8403 -197 8503 -181
rect 8561 -147 8661 -100
rect 8561 -181 8577 -147
rect 8645 -181 8661 -147
rect 8561 -197 8661 -181
rect 8719 -147 8819 -100
rect 8719 -181 8735 -147
rect 8803 -181 8819 -147
rect 8719 -197 8819 -181
rect 8877 -147 8977 -100
rect 8877 -181 8893 -147
rect 8961 -181 8977 -147
rect 8877 -197 8977 -181
rect 9035 -147 9135 -100
rect 9035 -181 9051 -147
rect 9119 -181 9135 -147
rect 9035 -197 9135 -181
rect 9193 -147 9293 -100
rect 9193 -181 9209 -147
rect 9277 -181 9293 -147
rect 9193 -197 9293 -181
rect 9351 -147 9451 -100
rect 9351 -181 9367 -147
rect 9435 -181 9451 -147
rect 9351 -197 9451 -181
rect 9509 -147 9609 -100
rect 9509 -181 9525 -147
rect 9593 -181 9609 -147
rect 9509 -197 9609 -181
rect 9667 -147 9767 -100
rect 9667 -181 9683 -147
rect 9751 -181 9767 -147
rect 9667 -197 9767 -181
rect 9825 -147 9925 -100
rect 9825 -181 9841 -147
rect 9909 -181 9925 -147
rect 9825 -197 9925 -181
rect 9983 -147 10083 -100
rect 9983 -181 9999 -147
rect 10067 -181 10083 -147
rect 9983 -197 10083 -181
rect 10141 -147 10241 -100
rect 10141 -181 10157 -147
rect 10225 -181 10241 -147
rect 10141 -197 10241 -181
rect 10299 -147 10399 -100
rect 10299 -181 10315 -147
rect 10383 -181 10399 -147
rect 10299 -197 10399 -181
rect 10457 -147 10557 -100
rect 10457 -181 10473 -147
rect 10541 -181 10557 -147
rect 10457 -197 10557 -181
rect 10615 -147 10715 -100
rect 10615 -181 10631 -147
rect 10699 -181 10715 -147
rect 10615 -197 10715 -181
rect 10773 -147 10873 -100
rect 10773 -181 10789 -147
rect 10857 -181 10873 -147
rect 10773 -197 10873 -181
rect 10931 -147 11031 -100
rect 10931 -181 10947 -147
rect 11015 -181 11031 -147
rect 10931 -197 11031 -181
rect 11089 -147 11189 -100
rect 11089 -181 11105 -147
rect 11173 -181 11189 -147
rect 11089 -197 11189 -181
rect 11247 -147 11347 -100
rect 11247 -181 11263 -147
rect 11331 -181 11347 -147
rect 11247 -197 11347 -181
rect 11405 -147 11505 -100
rect 11405 -181 11421 -147
rect 11489 -181 11505 -147
rect 11405 -197 11505 -181
rect 11563 -147 11663 -100
rect 11563 -181 11579 -147
rect 11647 -181 11663 -147
rect 11563 -197 11663 -181
rect 11721 -147 11821 -100
rect 11721 -181 11737 -147
rect 11805 -181 11821 -147
rect 11721 -197 11821 -181
rect 11879 -147 11979 -100
rect 11879 -181 11895 -147
rect 11963 -181 11979 -147
rect 11879 -197 11979 -181
rect 12037 -147 12137 -100
rect 12037 -181 12053 -147
rect 12121 -181 12137 -147
rect 12037 -197 12137 -181
rect 12195 -147 12295 -100
rect 12195 -181 12211 -147
rect 12279 -181 12295 -147
rect 12195 -197 12295 -181
rect 12353 -147 12453 -100
rect 12353 -181 12369 -147
rect 12437 -181 12453 -147
rect 12353 -197 12453 -181
rect 12511 -147 12611 -100
rect 12511 -181 12527 -147
rect 12595 -181 12611 -147
rect 12511 -197 12611 -181
rect 12669 -147 12769 -100
rect 12669 -181 12685 -147
rect 12753 -181 12769 -147
rect 12669 -197 12769 -181
rect 12827 -147 12927 -100
rect 12827 -181 12843 -147
rect 12911 -181 12927 -147
rect 12827 -197 12927 -181
rect 12985 -147 13085 -100
rect 12985 -181 13001 -147
rect 13069 -181 13085 -147
rect 12985 -197 13085 -181
rect 13143 -147 13243 -100
rect 13143 -181 13159 -147
rect 13227 -181 13243 -147
rect 13143 -197 13243 -181
rect 13301 -147 13401 -100
rect 13301 -181 13317 -147
rect 13385 -181 13401 -147
rect 13301 -197 13401 -181
rect 13459 -147 13559 -100
rect 13459 -181 13475 -147
rect 13543 -181 13559 -147
rect 13459 -197 13559 -181
rect 13617 -147 13717 -100
rect 13617 -181 13633 -147
rect 13701 -181 13717 -147
rect 13617 -197 13717 -181
rect 13775 -147 13875 -100
rect 13775 -181 13791 -147
rect 13859 -181 13875 -147
rect 13775 -197 13875 -181
rect 13933 -147 14033 -100
rect 13933 -181 13949 -147
rect 14017 -181 14033 -147
rect 13933 -197 14033 -181
rect 14091 -147 14191 -100
rect 14091 -181 14107 -147
rect 14175 -181 14191 -147
rect 14091 -197 14191 -181
rect 14249 -147 14349 -100
rect 14249 -181 14265 -147
rect 14333 -181 14349 -147
rect 14249 -197 14349 -181
rect 14407 -147 14507 -100
rect 14407 -181 14423 -147
rect 14491 -181 14507 -147
rect 14407 -197 14507 -181
rect 14565 -147 14665 -100
rect 14565 -181 14581 -147
rect 14649 -181 14665 -147
rect 14565 -197 14665 -181
rect 14723 -147 14823 -100
rect 14723 -181 14739 -147
rect 14807 -181 14823 -147
rect 14723 -197 14823 -181
rect 14881 -147 14981 -100
rect 14881 -181 14897 -147
rect 14965 -181 14981 -147
rect 14881 -197 14981 -181
rect 15039 -147 15139 -100
rect 15039 -181 15055 -147
rect 15123 -181 15139 -147
rect 15039 -197 15139 -181
rect 15197 -147 15297 -100
rect 15197 -181 15213 -147
rect 15281 -181 15297 -147
rect 15197 -197 15297 -181
rect 15355 -147 15455 -100
rect 15355 -181 15371 -147
rect 15439 -181 15455 -147
rect 15355 -197 15455 -181
rect 15513 -147 15613 -100
rect 15513 -181 15529 -147
rect 15597 -181 15613 -147
rect 15513 -197 15613 -181
rect 15671 -147 15771 -100
rect 15671 -181 15687 -147
rect 15755 -181 15771 -147
rect 15671 -197 15771 -181
<< polycont >>
rect -15755 147 -15687 181
rect -15597 147 -15529 181
rect -15439 147 -15371 181
rect -15281 147 -15213 181
rect -15123 147 -15055 181
rect -14965 147 -14897 181
rect -14807 147 -14739 181
rect -14649 147 -14581 181
rect -14491 147 -14423 181
rect -14333 147 -14265 181
rect -14175 147 -14107 181
rect -14017 147 -13949 181
rect -13859 147 -13791 181
rect -13701 147 -13633 181
rect -13543 147 -13475 181
rect -13385 147 -13317 181
rect -13227 147 -13159 181
rect -13069 147 -13001 181
rect -12911 147 -12843 181
rect -12753 147 -12685 181
rect -12595 147 -12527 181
rect -12437 147 -12369 181
rect -12279 147 -12211 181
rect -12121 147 -12053 181
rect -11963 147 -11895 181
rect -11805 147 -11737 181
rect -11647 147 -11579 181
rect -11489 147 -11421 181
rect -11331 147 -11263 181
rect -11173 147 -11105 181
rect -11015 147 -10947 181
rect -10857 147 -10789 181
rect -10699 147 -10631 181
rect -10541 147 -10473 181
rect -10383 147 -10315 181
rect -10225 147 -10157 181
rect -10067 147 -9999 181
rect -9909 147 -9841 181
rect -9751 147 -9683 181
rect -9593 147 -9525 181
rect -9435 147 -9367 181
rect -9277 147 -9209 181
rect -9119 147 -9051 181
rect -8961 147 -8893 181
rect -8803 147 -8735 181
rect -8645 147 -8577 181
rect -8487 147 -8419 181
rect -8329 147 -8261 181
rect -8171 147 -8103 181
rect -8013 147 -7945 181
rect -7855 147 -7787 181
rect -7697 147 -7629 181
rect -7539 147 -7471 181
rect -7381 147 -7313 181
rect -7223 147 -7155 181
rect -7065 147 -6997 181
rect -6907 147 -6839 181
rect -6749 147 -6681 181
rect -6591 147 -6523 181
rect -6433 147 -6365 181
rect -6275 147 -6207 181
rect -6117 147 -6049 181
rect -5959 147 -5891 181
rect -5801 147 -5733 181
rect -5643 147 -5575 181
rect -5485 147 -5417 181
rect -5327 147 -5259 181
rect -5169 147 -5101 181
rect -5011 147 -4943 181
rect -4853 147 -4785 181
rect -4695 147 -4627 181
rect -4537 147 -4469 181
rect -4379 147 -4311 181
rect -4221 147 -4153 181
rect -4063 147 -3995 181
rect -3905 147 -3837 181
rect -3747 147 -3679 181
rect -3589 147 -3521 181
rect -3431 147 -3363 181
rect -3273 147 -3205 181
rect -3115 147 -3047 181
rect -2957 147 -2889 181
rect -2799 147 -2731 181
rect -2641 147 -2573 181
rect -2483 147 -2415 181
rect -2325 147 -2257 181
rect -2167 147 -2099 181
rect -2009 147 -1941 181
rect -1851 147 -1783 181
rect -1693 147 -1625 181
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect 1625 147 1693 181
rect 1783 147 1851 181
rect 1941 147 2009 181
rect 2099 147 2167 181
rect 2257 147 2325 181
rect 2415 147 2483 181
rect 2573 147 2641 181
rect 2731 147 2799 181
rect 2889 147 2957 181
rect 3047 147 3115 181
rect 3205 147 3273 181
rect 3363 147 3431 181
rect 3521 147 3589 181
rect 3679 147 3747 181
rect 3837 147 3905 181
rect 3995 147 4063 181
rect 4153 147 4221 181
rect 4311 147 4379 181
rect 4469 147 4537 181
rect 4627 147 4695 181
rect 4785 147 4853 181
rect 4943 147 5011 181
rect 5101 147 5169 181
rect 5259 147 5327 181
rect 5417 147 5485 181
rect 5575 147 5643 181
rect 5733 147 5801 181
rect 5891 147 5959 181
rect 6049 147 6117 181
rect 6207 147 6275 181
rect 6365 147 6433 181
rect 6523 147 6591 181
rect 6681 147 6749 181
rect 6839 147 6907 181
rect 6997 147 7065 181
rect 7155 147 7223 181
rect 7313 147 7381 181
rect 7471 147 7539 181
rect 7629 147 7697 181
rect 7787 147 7855 181
rect 7945 147 8013 181
rect 8103 147 8171 181
rect 8261 147 8329 181
rect 8419 147 8487 181
rect 8577 147 8645 181
rect 8735 147 8803 181
rect 8893 147 8961 181
rect 9051 147 9119 181
rect 9209 147 9277 181
rect 9367 147 9435 181
rect 9525 147 9593 181
rect 9683 147 9751 181
rect 9841 147 9909 181
rect 9999 147 10067 181
rect 10157 147 10225 181
rect 10315 147 10383 181
rect 10473 147 10541 181
rect 10631 147 10699 181
rect 10789 147 10857 181
rect 10947 147 11015 181
rect 11105 147 11173 181
rect 11263 147 11331 181
rect 11421 147 11489 181
rect 11579 147 11647 181
rect 11737 147 11805 181
rect 11895 147 11963 181
rect 12053 147 12121 181
rect 12211 147 12279 181
rect 12369 147 12437 181
rect 12527 147 12595 181
rect 12685 147 12753 181
rect 12843 147 12911 181
rect 13001 147 13069 181
rect 13159 147 13227 181
rect 13317 147 13385 181
rect 13475 147 13543 181
rect 13633 147 13701 181
rect 13791 147 13859 181
rect 13949 147 14017 181
rect 14107 147 14175 181
rect 14265 147 14333 181
rect 14423 147 14491 181
rect 14581 147 14649 181
rect 14739 147 14807 181
rect 14897 147 14965 181
rect 15055 147 15123 181
rect 15213 147 15281 181
rect 15371 147 15439 181
rect 15529 147 15597 181
rect 15687 147 15755 181
rect -15755 -181 -15687 -147
rect -15597 -181 -15529 -147
rect -15439 -181 -15371 -147
rect -15281 -181 -15213 -147
rect -15123 -181 -15055 -147
rect -14965 -181 -14897 -147
rect -14807 -181 -14739 -147
rect -14649 -181 -14581 -147
rect -14491 -181 -14423 -147
rect -14333 -181 -14265 -147
rect -14175 -181 -14107 -147
rect -14017 -181 -13949 -147
rect -13859 -181 -13791 -147
rect -13701 -181 -13633 -147
rect -13543 -181 -13475 -147
rect -13385 -181 -13317 -147
rect -13227 -181 -13159 -147
rect -13069 -181 -13001 -147
rect -12911 -181 -12843 -147
rect -12753 -181 -12685 -147
rect -12595 -181 -12527 -147
rect -12437 -181 -12369 -147
rect -12279 -181 -12211 -147
rect -12121 -181 -12053 -147
rect -11963 -181 -11895 -147
rect -11805 -181 -11737 -147
rect -11647 -181 -11579 -147
rect -11489 -181 -11421 -147
rect -11331 -181 -11263 -147
rect -11173 -181 -11105 -147
rect -11015 -181 -10947 -147
rect -10857 -181 -10789 -147
rect -10699 -181 -10631 -147
rect -10541 -181 -10473 -147
rect -10383 -181 -10315 -147
rect -10225 -181 -10157 -147
rect -10067 -181 -9999 -147
rect -9909 -181 -9841 -147
rect -9751 -181 -9683 -147
rect -9593 -181 -9525 -147
rect -9435 -181 -9367 -147
rect -9277 -181 -9209 -147
rect -9119 -181 -9051 -147
rect -8961 -181 -8893 -147
rect -8803 -181 -8735 -147
rect -8645 -181 -8577 -147
rect -8487 -181 -8419 -147
rect -8329 -181 -8261 -147
rect -8171 -181 -8103 -147
rect -8013 -181 -7945 -147
rect -7855 -181 -7787 -147
rect -7697 -181 -7629 -147
rect -7539 -181 -7471 -147
rect -7381 -181 -7313 -147
rect -7223 -181 -7155 -147
rect -7065 -181 -6997 -147
rect -6907 -181 -6839 -147
rect -6749 -181 -6681 -147
rect -6591 -181 -6523 -147
rect -6433 -181 -6365 -147
rect -6275 -181 -6207 -147
rect -6117 -181 -6049 -147
rect -5959 -181 -5891 -147
rect -5801 -181 -5733 -147
rect -5643 -181 -5575 -147
rect -5485 -181 -5417 -147
rect -5327 -181 -5259 -147
rect -5169 -181 -5101 -147
rect -5011 -181 -4943 -147
rect -4853 -181 -4785 -147
rect -4695 -181 -4627 -147
rect -4537 -181 -4469 -147
rect -4379 -181 -4311 -147
rect -4221 -181 -4153 -147
rect -4063 -181 -3995 -147
rect -3905 -181 -3837 -147
rect -3747 -181 -3679 -147
rect -3589 -181 -3521 -147
rect -3431 -181 -3363 -147
rect -3273 -181 -3205 -147
rect -3115 -181 -3047 -147
rect -2957 -181 -2889 -147
rect -2799 -181 -2731 -147
rect -2641 -181 -2573 -147
rect -2483 -181 -2415 -147
rect -2325 -181 -2257 -147
rect -2167 -181 -2099 -147
rect -2009 -181 -1941 -147
rect -1851 -181 -1783 -147
rect -1693 -181 -1625 -147
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
rect 1625 -181 1693 -147
rect 1783 -181 1851 -147
rect 1941 -181 2009 -147
rect 2099 -181 2167 -147
rect 2257 -181 2325 -147
rect 2415 -181 2483 -147
rect 2573 -181 2641 -147
rect 2731 -181 2799 -147
rect 2889 -181 2957 -147
rect 3047 -181 3115 -147
rect 3205 -181 3273 -147
rect 3363 -181 3431 -147
rect 3521 -181 3589 -147
rect 3679 -181 3747 -147
rect 3837 -181 3905 -147
rect 3995 -181 4063 -147
rect 4153 -181 4221 -147
rect 4311 -181 4379 -147
rect 4469 -181 4537 -147
rect 4627 -181 4695 -147
rect 4785 -181 4853 -147
rect 4943 -181 5011 -147
rect 5101 -181 5169 -147
rect 5259 -181 5327 -147
rect 5417 -181 5485 -147
rect 5575 -181 5643 -147
rect 5733 -181 5801 -147
rect 5891 -181 5959 -147
rect 6049 -181 6117 -147
rect 6207 -181 6275 -147
rect 6365 -181 6433 -147
rect 6523 -181 6591 -147
rect 6681 -181 6749 -147
rect 6839 -181 6907 -147
rect 6997 -181 7065 -147
rect 7155 -181 7223 -147
rect 7313 -181 7381 -147
rect 7471 -181 7539 -147
rect 7629 -181 7697 -147
rect 7787 -181 7855 -147
rect 7945 -181 8013 -147
rect 8103 -181 8171 -147
rect 8261 -181 8329 -147
rect 8419 -181 8487 -147
rect 8577 -181 8645 -147
rect 8735 -181 8803 -147
rect 8893 -181 8961 -147
rect 9051 -181 9119 -147
rect 9209 -181 9277 -147
rect 9367 -181 9435 -147
rect 9525 -181 9593 -147
rect 9683 -181 9751 -147
rect 9841 -181 9909 -147
rect 9999 -181 10067 -147
rect 10157 -181 10225 -147
rect 10315 -181 10383 -147
rect 10473 -181 10541 -147
rect 10631 -181 10699 -147
rect 10789 -181 10857 -147
rect 10947 -181 11015 -147
rect 11105 -181 11173 -147
rect 11263 -181 11331 -147
rect 11421 -181 11489 -147
rect 11579 -181 11647 -147
rect 11737 -181 11805 -147
rect 11895 -181 11963 -147
rect 12053 -181 12121 -147
rect 12211 -181 12279 -147
rect 12369 -181 12437 -147
rect 12527 -181 12595 -147
rect 12685 -181 12753 -147
rect 12843 -181 12911 -147
rect 13001 -181 13069 -147
rect 13159 -181 13227 -147
rect 13317 -181 13385 -147
rect 13475 -181 13543 -147
rect 13633 -181 13701 -147
rect 13791 -181 13859 -147
rect 13949 -181 14017 -147
rect 14107 -181 14175 -147
rect 14265 -181 14333 -147
rect 14423 -181 14491 -147
rect 14581 -181 14649 -147
rect 14739 -181 14807 -147
rect 14897 -181 14965 -147
rect 15055 -181 15123 -147
rect 15213 -181 15281 -147
rect 15371 -181 15439 -147
rect 15529 -181 15597 -147
rect 15687 -181 15755 -147
<< locali >>
rect -15951 285 -15855 319
rect 15855 285 15951 319
rect -15951 223 -15917 285
rect 15917 223 15951 285
rect -15771 147 -15755 181
rect -15687 147 -15671 181
rect -15613 147 -15597 181
rect -15529 147 -15513 181
rect -15455 147 -15439 181
rect -15371 147 -15355 181
rect -15297 147 -15281 181
rect -15213 147 -15197 181
rect -15139 147 -15123 181
rect -15055 147 -15039 181
rect -14981 147 -14965 181
rect -14897 147 -14881 181
rect -14823 147 -14807 181
rect -14739 147 -14723 181
rect -14665 147 -14649 181
rect -14581 147 -14565 181
rect -14507 147 -14491 181
rect -14423 147 -14407 181
rect -14349 147 -14333 181
rect -14265 147 -14249 181
rect -14191 147 -14175 181
rect -14107 147 -14091 181
rect -14033 147 -14017 181
rect -13949 147 -13933 181
rect -13875 147 -13859 181
rect -13791 147 -13775 181
rect -13717 147 -13701 181
rect -13633 147 -13617 181
rect -13559 147 -13543 181
rect -13475 147 -13459 181
rect -13401 147 -13385 181
rect -13317 147 -13301 181
rect -13243 147 -13227 181
rect -13159 147 -13143 181
rect -13085 147 -13069 181
rect -13001 147 -12985 181
rect -12927 147 -12911 181
rect -12843 147 -12827 181
rect -12769 147 -12753 181
rect -12685 147 -12669 181
rect -12611 147 -12595 181
rect -12527 147 -12511 181
rect -12453 147 -12437 181
rect -12369 147 -12353 181
rect -12295 147 -12279 181
rect -12211 147 -12195 181
rect -12137 147 -12121 181
rect -12053 147 -12037 181
rect -11979 147 -11963 181
rect -11895 147 -11879 181
rect -11821 147 -11805 181
rect -11737 147 -11721 181
rect -11663 147 -11647 181
rect -11579 147 -11563 181
rect -11505 147 -11489 181
rect -11421 147 -11405 181
rect -11347 147 -11331 181
rect -11263 147 -11247 181
rect -11189 147 -11173 181
rect -11105 147 -11089 181
rect -11031 147 -11015 181
rect -10947 147 -10931 181
rect -10873 147 -10857 181
rect -10789 147 -10773 181
rect -10715 147 -10699 181
rect -10631 147 -10615 181
rect -10557 147 -10541 181
rect -10473 147 -10457 181
rect -10399 147 -10383 181
rect -10315 147 -10299 181
rect -10241 147 -10225 181
rect -10157 147 -10141 181
rect -10083 147 -10067 181
rect -9999 147 -9983 181
rect -9925 147 -9909 181
rect -9841 147 -9825 181
rect -9767 147 -9751 181
rect -9683 147 -9667 181
rect -9609 147 -9593 181
rect -9525 147 -9509 181
rect -9451 147 -9435 181
rect -9367 147 -9351 181
rect -9293 147 -9277 181
rect -9209 147 -9193 181
rect -9135 147 -9119 181
rect -9051 147 -9035 181
rect -8977 147 -8961 181
rect -8893 147 -8877 181
rect -8819 147 -8803 181
rect -8735 147 -8719 181
rect -8661 147 -8645 181
rect -8577 147 -8561 181
rect -8503 147 -8487 181
rect -8419 147 -8403 181
rect -8345 147 -8329 181
rect -8261 147 -8245 181
rect -8187 147 -8171 181
rect -8103 147 -8087 181
rect -8029 147 -8013 181
rect -7945 147 -7929 181
rect -7871 147 -7855 181
rect -7787 147 -7771 181
rect -7713 147 -7697 181
rect -7629 147 -7613 181
rect -7555 147 -7539 181
rect -7471 147 -7455 181
rect -7397 147 -7381 181
rect -7313 147 -7297 181
rect -7239 147 -7223 181
rect -7155 147 -7139 181
rect -7081 147 -7065 181
rect -6997 147 -6981 181
rect -6923 147 -6907 181
rect -6839 147 -6823 181
rect -6765 147 -6749 181
rect -6681 147 -6665 181
rect -6607 147 -6591 181
rect -6523 147 -6507 181
rect -6449 147 -6433 181
rect -6365 147 -6349 181
rect -6291 147 -6275 181
rect -6207 147 -6191 181
rect -6133 147 -6117 181
rect -6049 147 -6033 181
rect -5975 147 -5959 181
rect -5891 147 -5875 181
rect -5817 147 -5801 181
rect -5733 147 -5717 181
rect -5659 147 -5643 181
rect -5575 147 -5559 181
rect -5501 147 -5485 181
rect -5417 147 -5401 181
rect -5343 147 -5327 181
rect -5259 147 -5243 181
rect -5185 147 -5169 181
rect -5101 147 -5085 181
rect -5027 147 -5011 181
rect -4943 147 -4927 181
rect -4869 147 -4853 181
rect -4785 147 -4769 181
rect -4711 147 -4695 181
rect -4627 147 -4611 181
rect -4553 147 -4537 181
rect -4469 147 -4453 181
rect -4395 147 -4379 181
rect -4311 147 -4295 181
rect -4237 147 -4221 181
rect -4153 147 -4137 181
rect -4079 147 -4063 181
rect -3995 147 -3979 181
rect -3921 147 -3905 181
rect -3837 147 -3821 181
rect -3763 147 -3747 181
rect -3679 147 -3663 181
rect -3605 147 -3589 181
rect -3521 147 -3505 181
rect -3447 147 -3431 181
rect -3363 147 -3347 181
rect -3289 147 -3273 181
rect -3205 147 -3189 181
rect -3131 147 -3115 181
rect -3047 147 -3031 181
rect -2973 147 -2957 181
rect -2889 147 -2873 181
rect -2815 147 -2799 181
rect -2731 147 -2715 181
rect -2657 147 -2641 181
rect -2573 147 -2557 181
rect -2499 147 -2483 181
rect -2415 147 -2399 181
rect -2341 147 -2325 181
rect -2257 147 -2241 181
rect -2183 147 -2167 181
rect -2099 147 -2083 181
rect -2025 147 -2009 181
rect -1941 147 -1925 181
rect -1867 147 -1851 181
rect -1783 147 -1767 181
rect -1709 147 -1693 181
rect -1625 147 -1609 181
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -919 147 -903 181
rect -835 147 -819 181
rect -761 147 -745 181
rect -677 147 -661 181
rect -603 147 -587 181
rect -519 147 -503 181
rect -445 147 -429 181
rect -361 147 -345 181
rect -287 147 -271 181
rect -203 147 -187 181
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect 187 147 203 181
rect 271 147 287 181
rect 345 147 361 181
rect 429 147 445 181
rect 503 147 519 181
rect 587 147 603 181
rect 661 147 677 181
rect 745 147 761 181
rect 819 147 835 181
rect 903 147 919 181
rect 977 147 993 181
rect 1061 147 1077 181
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1451 147 1467 181
rect 1535 147 1551 181
rect 1609 147 1625 181
rect 1693 147 1709 181
rect 1767 147 1783 181
rect 1851 147 1867 181
rect 1925 147 1941 181
rect 2009 147 2025 181
rect 2083 147 2099 181
rect 2167 147 2183 181
rect 2241 147 2257 181
rect 2325 147 2341 181
rect 2399 147 2415 181
rect 2483 147 2499 181
rect 2557 147 2573 181
rect 2641 147 2657 181
rect 2715 147 2731 181
rect 2799 147 2815 181
rect 2873 147 2889 181
rect 2957 147 2973 181
rect 3031 147 3047 181
rect 3115 147 3131 181
rect 3189 147 3205 181
rect 3273 147 3289 181
rect 3347 147 3363 181
rect 3431 147 3447 181
rect 3505 147 3521 181
rect 3589 147 3605 181
rect 3663 147 3679 181
rect 3747 147 3763 181
rect 3821 147 3837 181
rect 3905 147 3921 181
rect 3979 147 3995 181
rect 4063 147 4079 181
rect 4137 147 4153 181
rect 4221 147 4237 181
rect 4295 147 4311 181
rect 4379 147 4395 181
rect 4453 147 4469 181
rect 4537 147 4553 181
rect 4611 147 4627 181
rect 4695 147 4711 181
rect 4769 147 4785 181
rect 4853 147 4869 181
rect 4927 147 4943 181
rect 5011 147 5027 181
rect 5085 147 5101 181
rect 5169 147 5185 181
rect 5243 147 5259 181
rect 5327 147 5343 181
rect 5401 147 5417 181
rect 5485 147 5501 181
rect 5559 147 5575 181
rect 5643 147 5659 181
rect 5717 147 5733 181
rect 5801 147 5817 181
rect 5875 147 5891 181
rect 5959 147 5975 181
rect 6033 147 6049 181
rect 6117 147 6133 181
rect 6191 147 6207 181
rect 6275 147 6291 181
rect 6349 147 6365 181
rect 6433 147 6449 181
rect 6507 147 6523 181
rect 6591 147 6607 181
rect 6665 147 6681 181
rect 6749 147 6765 181
rect 6823 147 6839 181
rect 6907 147 6923 181
rect 6981 147 6997 181
rect 7065 147 7081 181
rect 7139 147 7155 181
rect 7223 147 7239 181
rect 7297 147 7313 181
rect 7381 147 7397 181
rect 7455 147 7471 181
rect 7539 147 7555 181
rect 7613 147 7629 181
rect 7697 147 7713 181
rect 7771 147 7787 181
rect 7855 147 7871 181
rect 7929 147 7945 181
rect 8013 147 8029 181
rect 8087 147 8103 181
rect 8171 147 8187 181
rect 8245 147 8261 181
rect 8329 147 8345 181
rect 8403 147 8419 181
rect 8487 147 8503 181
rect 8561 147 8577 181
rect 8645 147 8661 181
rect 8719 147 8735 181
rect 8803 147 8819 181
rect 8877 147 8893 181
rect 8961 147 8977 181
rect 9035 147 9051 181
rect 9119 147 9135 181
rect 9193 147 9209 181
rect 9277 147 9293 181
rect 9351 147 9367 181
rect 9435 147 9451 181
rect 9509 147 9525 181
rect 9593 147 9609 181
rect 9667 147 9683 181
rect 9751 147 9767 181
rect 9825 147 9841 181
rect 9909 147 9925 181
rect 9983 147 9999 181
rect 10067 147 10083 181
rect 10141 147 10157 181
rect 10225 147 10241 181
rect 10299 147 10315 181
rect 10383 147 10399 181
rect 10457 147 10473 181
rect 10541 147 10557 181
rect 10615 147 10631 181
rect 10699 147 10715 181
rect 10773 147 10789 181
rect 10857 147 10873 181
rect 10931 147 10947 181
rect 11015 147 11031 181
rect 11089 147 11105 181
rect 11173 147 11189 181
rect 11247 147 11263 181
rect 11331 147 11347 181
rect 11405 147 11421 181
rect 11489 147 11505 181
rect 11563 147 11579 181
rect 11647 147 11663 181
rect 11721 147 11737 181
rect 11805 147 11821 181
rect 11879 147 11895 181
rect 11963 147 11979 181
rect 12037 147 12053 181
rect 12121 147 12137 181
rect 12195 147 12211 181
rect 12279 147 12295 181
rect 12353 147 12369 181
rect 12437 147 12453 181
rect 12511 147 12527 181
rect 12595 147 12611 181
rect 12669 147 12685 181
rect 12753 147 12769 181
rect 12827 147 12843 181
rect 12911 147 12927 181
rect 12985 147 13001 181
rect 13069 147 13085 181
rect 13143 147 13159 181
rect 13227 147 13243 181
rect 13301 147 13317 181
rect 13385 147 13401 181
rect 13459 147 13475 181
rect 13543 147 13559 181
rect 13617 147 13633 181
rect 13701 147 13717 181
rect 13775 147 13791 181
rect 13859 147 13875 181
rect 13933 147 13949 181
rect 14017 147 14033 181
rect 14091 147 14107 181
rect 14175 147 14191 181
rect 14249 147 14265 181
rect 14333 147 14349 181
rect 14407 147 14423 181
rect 14491 147 14507 181
rect 14565 147 14581 181
rect 14649 147 14665 181
rect 14723 147 14739 181
rect 14807 147 14823 181
rect 14881 147 14897 181
rect 14965 147 14981 181
rect 15039 147 15055 181
rect 15123 147 15139 181
rect 15197 147 15213 181
rect 15281 147 15297 181
rect 15355 147 15371 181
rect 15439 147 15455 181
rect 15513 147 15529 181
rect 15597 147 15613 181
rect 15671 147 15687 181
rect 15755 147 15771 181
rect -15817 88 -15783 104
rect -15817 -104 -15783 -88
rect -15659 88 -15625 104
rect -15659 -104 -15625 -88
rect -15501 88 -15467 104
rect -15501 -104 -15467 -88
rect -15343 88 -15309 104
rect -15343 -104 -15309 -88
rect -15185 88 -15151 104
rect -15185 -104 -15151 -88
rect -15027 88 -14993 104
rect -15027 -104 -14993 -88
rect -14869 88 -14835 104
rect -14869 -104 -14835 -88
rect -14711 88 -14677 104
rect -14711 -104 -14677 -88
rect -14553 88 -14519 104
rect -14553 -104 -14519 -88
rect -14395 88 -14361 104
rect -14395 -104 -14361 -88
rect -14237 88 -14203 104
rect -14237 -104 -14203 -88
rect -14079 88 -14045 104
rect -14079 -104 -14045 -88
rect -13921 88 -13887 104
rect -13921 -104 -13887 -88
rect -13763 88 -13729 104
rect -13763 -104 -13729 -88
rect -13605 88 -13571 104
rect -13605 -104 -13571 -88
rect -13447 88 -13413 104
rect -13447 -104 -13413 -88
rect -13289 88 -13255 104
rect -13289 -104 -13255 -88
rect -13131 88 -13097 104
rect -13131 -104 -13097 -88
rect -12973 88 -12939 104
rect -12973 -104 -12939 -88
rect -12815 88 -12781 104
rect -12815 -104 -12781 -88
rect -12657 88 -12623 104
rect -12657 -104 -12623 -88
rect -12499 88 -12465 104
rect -12499 -104 -12465 -88
rect -12341 88 -12307 104
rect -12341 -104 -12307 -88
rect -12183 88 -12149 104
rect -12183 -104 -12149 -88
rect -12025 88 -11991 104
rect -12025 -104 -11991 -88
rect -11867 88 -11833 104
rect -11867 -104 -11833 -88
rect -11709 88 -11675 104
rect -11709 -104 -11675 -88
rect -11551 88 -11517 104
rect -11551 -104 -11517 -88
rect -11393 88 -11359 104
rect -11393 -104 -11359 -88
rect -11235 88 -11201 104
rect -11235 -104 -11201 -88
rect -11077 88 -11043 104
rect -11077 -104 -11043 -88
rect -10919 88 -10885 104
rect -10919 -104 -10885 -88
rect -10761 88 -10727 104
rect -10761 -104 -10727 -88
rect -10603 88 -10569 104
rect -10603 -104 -10569 -88
rect -10445 88 -10411 104
rect -10445 -104 -10411 -88
rect -10287 88 -10253 104
rect -10287 -104 -10253 -88
rect -10129 88 -10095 104
rect -10129 -104 -10095 -88
rect -9971 88 -9937 104
rect -9971 -104 -9937 -88
rect -9813 88 -9779 104
rect -9813 -104 -9779 -88
rect -9655 88 -9621 104
rect -9655 -104 -9621 -88
rect -9497 88 -9463 104
rect -9497 -104 -9463 -88
rect -9339 88 -9305 104
rect -9339 -104 -9305 -88
rect -9181 88 -9147 104
rect -9181 -104 -9147 -88
rect -9023 88 -8989 104
rect -9023 -104 -8989 -88
rect -8865 88 -8831 104
rect -8865 -104 -8831 -88
rect -8707 88 -8673 104
rect -8707 -104 -8673 -88
rect -8549 88 -8515 104
rect -8549 -104 -8515 -88
rect -8391 88 -8357 104
rect -8391 -104 -8357 -88
rect -8233 88 -8199 104
rect -8233 -104 -8199 -88
rect -8075 88 -8041 104
rect -8075 -104 -8041 -88
rect -7917 88 -7883 104
rect -7917 -104 -7883 -88
rect -7759 88 -7725 104
rect -7759 -104 -7725 -88
rect -7601 88 -7567 104
rect -7601 -104 -7567 -88
rect -7443 88 -7409 104
rect -7443 -104 -7409 -88
rect -7285 88 -7251 104
rect -7285 -104 -7251 -88
rect -7127 88 -7093 104
rect -7127 -104 -7093 -88
rect -6969 88 -6935 104
rect -6969 -104 -6935 -88
rect -6811 88 -6777 104
rect -6811 -104 -6777 -88
rect -6653 88 -6619 104
rect -6653 -104 -6619 -88
rect -6495 88 -6461 104
rect -6495 -104 -6461 -88
rect -6337 88 -6303 104
rect -6337 -104 -6303 -88
rect -6179 88 -6145 104
rect -6179 -104 -6145 -88
rect -6021 88 -5987 104
rect -6021 -104 -5987 -88
rect -5863 88 -5829 104
rect -5863 -104 -5829 -88
rect -5705 88 -5671 104
rect -5705 -104 -5671 -88
rect -5547 88 -5513 104
rect -5547 -104 -5513 -88
rect -5389 88 -5355 104
rect -5389 -104 -5355 -88
rect -5231 88 -5197 104
rect -5231 -104 -5197 -88
rect -5073 88 -5039 104
rect -5073 -104 -5039 -88
rect -4915 88 -4881 104
rect -4915 -104 -4881 -88
rect -4757 88 -4723 104
rect -4757 -104 -4723 -88
rect -4599 88 -4565 104
rect -4599 -104 -4565 -88
rect -4441 88 -4407 104
rect -4441 -104 -4407 -88
rect -4283 88 -4249 104
rect -4283 -104 -4249 -88
rect -4125 88 -4091 104
rect -4125 -104 -4091 -88
rect -3967 88 -3933 104
rect -3967 -104 -3933 -88
rect -3809 88 -3775 104
rect -3809 -104 -3775 -88
rect -3651 88 -3617 104
rect -3651 -104 -3617 -88
rect -3493 88 -3459 104
rect -3493 -104 -3459 -88
rect -3335 88 -3301 104
rect -3335 -104 -3301 -88
rect -3177 88 -3143 104
rect -3177 -104 -3143 -88
rect -3019 88 -2985 104
rect -3019 -104 -2985 -88
rect -2861 88 -2827 104
rect -2861 -104 -2827 -88
rect -2703 88 -2669 104
rect -2703 -104 -2669 -88
rect -2545 88 -2511 104
rect -2545 -104 -2511 -88
rect -2387 88 -2353 104
rect -2387 -104 -2353 -88
rect -2229 88 -2195 104
rect -2229 -104 -2195 -88
rect -2071 88 -2037 104
rect -2071 -104 -2037 -88
rect -1913 88 -1879 104
rect -1913 -104 -1879 -88
rect -1755 88 -1721 104
rect -1755 -104 -1721 -88
rect -1597 88 -1563 104
rect -1597 -104 -1563 -88
rect -1439 88 -1405 104
rect -1439 -104 -1405 -88
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect 1405 88 1439 104
rect 1405 -104 1439 -88
rect 1563 88 1597 104
rect 1563 -104 1597 -88
rect 1721 88 1755 104
rect 1721 -104 1755 -88
rect 1879 88 1913 104
rect 1879 -104 1913 -88
rect 2037 88 2071 104
rect 2037 -104 2071 -88
rect 2195 88 2229 104
rect 2195 -104 2229 -88
rect 2353 88 2387 104
rect 2353 -104 2387 -88
rect 2511 88 2545 104
rect 2511 -104 2545 -88
rect 2669 88 2703 104
rect 2669 -104 2703 -88
rect 2827 88 2861 104
rect 2827 -104 2861 -88
rect 2985 88 3019 104
rect 2985 -104 3019 -88
rect 3143 88 3177 104
rect 3143 -104 3177 -88
rect 3301 88 3335 104
rect 3301 -104 3335 -88
rect 3459 88 3493 104
rect 3459 -104 3493 -88
rect 3617 88 3651 104
rect 3617 -104 3651 -88
rect 3775 88 3809 104
rect 3775 -104 3809 -88
rect 3933 88 3967 104
rect 3933 -104 3967 -88
rect 4091 88 4125 104
rect 4091 -104 4125 -88
rect 4249 88 4283 104
rect 4249 -104 4283 -88
rect 4407 88 4441 104
rect 4407 -104 4441 -88
rect 4565 88 4599 104
rect 4565 -104 4599 -88
rect 4723 88 4757 104
rect 4723 -104 4757 -88
rect 4881 88 4915 104
rect 4881 -104 4915 -88
rect 5039 88 5073 104
rect 5039 -104 5073 -88
rect 5197 88 5231 104
rect 5197 -104 5231 -88
rect 5355 88 5389 104
rect 5355 -104 5389 -88
rect 5513 88 5547 104
rect 5513 -104 5547 -88
rect 5671 88 5705 104
rect 5671 -104 5705 -88
rect 5829 88 5863 104
rect 5829 -104 5863 -88
rect 5987 88 6021 104
rect 5987 -104 6021 -88
rect 6145 88 6179 104
rect 6145 -104 6179 -88
rect 6303 88 6337 104
rect 6303 -104 6337 -88
rect 6461 88 6495 104
rect 6461 -104 6495 -88
rect 6619 88 6653 104
rect 6619 -104 6653 -88
rect 6777 88 6811 104
rect 6777 -104 6811 -88
rect 6935 88 6969 104
rect 6935 -104 6969 -88
rect 7093 88 7127 104
rect 7093 -104 7127 -88
rect 7251 88 7285 104
rect 7251 -104 7285 -88
rect 7409 88 7443 104
rect 7409 -104 7443 -88
rect 7567 88 7601 104
rect 7567 -104 7601 -88
rect 7725 88 7759 104
rect 7725 -104 7759 -88
rect 7883 88 7917 104
rect 7883 -104 7917 -88
rect 8041 88 8075 104
rect 8041 -104 8075 -88
rect 8199 88 8233 104
rect 8199 -104 8233 -88
rect 8357 88 8391 104
rect 8357 -104 8391 -88
rect 8515 88 8549 104
rect 8515 -104 8549 -88
rect 8673 88 8707 104
rect 8673 -104 8707 -88
rect 8831 88 8865 104
rect 8831 -104 8865 -88
rect 8989 88 9023 104
rect 8989 -104 9023 -88
rect 9147 88 9181 104
rect 9147 -104 9181 -88
rect 9305 88 9339 104
rect 9305 -104 9339 -88
rect 9463 88 9497 104
rect 9463 -104 9497 -88
rect 9621 88 9655 104
rect 9621 -104 9655 -88
rect 9779 88 9813 104
rect 9779 -104 9813 -88
rect 9937 88 9971 104
rect 9937 -104 9971 -88
rect 10095 88 10129 104
rect 10095 -104 10129 -88
rect 10253 88 10287 104
rect 10253 -104 10287 -88
rect 10411 88 10445 104
rect 10411 -104 10445 -88
rect 10569 88 10603 104
rect 10569 -104 10603 -88
rect 10727 88 10761 104
rect 10727 -104 10761 -88
rect 10885 88 10919 104
rect 10885 -104 10919 -88
rect 11043 88 11077 104
rect 11043 -104 11077 -88
rect 11201 88 11235 104
rect 11201 -104 11235 -88
rect 11359 88 11393 104
rect 11359 -104 11393 -88
rect 11517 88 11551 104
rect 11517 -104 11551 -88
rect 11675 88 11709 104
rect 11675 -104 11709 -88
rect 11833 88 11867 104
rect 11833 -104 11867 -88
rect 11991 88 12025 104
rect 11991 -104 12025 -88
rect 12149 88 12183 104
rect 12149 -104 12183 -88
rect 12307 88 12341 104
rect 12307 -104 12341 -88
rect 12465 88 12499 104
rect 12465 -104 12499 -88
rect 12623 88 12657 104
rect 12623 -104 12657 -88
rect 12781 88 12815 104
rect 12781 -104 12815 -88
rect 12939 88 12973 104
rect 12939 -104 12973 -88
rect 13097 88 13131 104
rect 13097 -104 13131 -88
rect 13255 88 13289 104
rect 13255 -104 13289 -88
rect 13413 88 13447 104
rect 13413 -104 13447 -88
rect 13571 88 13605 104
rect 13571 -104 13605 -88
rect 13729 88 13763 104
rect 13729 -104 13763 -88
rect 13887 88 13921 104
rect 13887 -104 13921 -88
rect 14045 88 14079 104
rect 14045 -104 14079 -88
rect 14203 88 14237 104
rect 14203 -104 14237 -88
rect 14361 88 14395 104
rect 14361 -104 14395 -88
rect 14519 88 14553 104
rect 14519 -104 14553 -88
rect 14677 88 14711 104
rect 14677 -104 14711 -88
rect 14835 88 14869 104
rect 14835 -104 14869 -88
rect 14993 88 15027 104
rect 14993 -104 15027 -88
rect 15151 88 15185 104
rect 15151 -104 15185 -88
rect 15309 88 15343 104
rect 15309 -104 15343 -88
rect 15467 88 15501 104
rect 15467 -104 15501 -88
rect 15625 88 15659 104
rect 15625 -104 15659 -88
rect 15783 88 15817 104
rect 15783 -104 15817 -88
rect -15771 -181 -15755 -147
rect -15687 -181 -15671 -147
rect -15613 -181 -15597 -147
rect -15529 -181 -15513 -147
rect -15455 -181 -15439 -147
rect -15371 -181 -15355 -147
rect -15297 -181 -15281 -147
rect -15213 -181 -15197 -147
rect -15139 -181 -15123 -147
rect -15055 -181 -15039 -147
rect -14981 -181 -14965 -147
rect -14897 -181 -14881 -147
rect -14823 -181 -14807 -147
rect -14739 -181 -14723 -147
rect -14665 -181 -14649 -147
rect -14581 -181 -14565 -147
rect -14507 -181 -14491 -147
rect -14423 -181 -14407 -147
rect -14349 -181 -14333 -147
rect -14265 -181 -14249 -147
rect -14191 -181 -14175 -147
rect -14107 -181 -14091 -147
rect -14033 -181 -14017 -147
rect -13949 -181 -13933 -147
rect -13875 -181 -13859 -147
rect -13791 -181 -13775 -147
rect -13717 -181 -13701 -147
rect -13633 -181 -13617 -147
rect -13559 -181 -13543 -147
rect -13475 -181 -13459 -147
rect -13401 -181 -13385 -147
rect -13317 -181 -13301 -147
rect -13243 -181 -13227 -147
rect -13159 -181 -13143 -147
rect -13085 -181 -13069 -147
rect -13001 -181 -12985 -147
rect -12927 -181 -12911 -147
rect -12843 -181 -12827 -147
rect -12769 -181 -12753 -147
rect -12685 -181 -12669 -147
rect -12611 -181 -12595 -147
rect -12527 -181 -12511 -147
rect -12453 -181 -12437 -147
rect -12369 -181 -12353 -147
rect -12295 -181 -12279 -147
rect -12211 -181 -12195 -147
rect -12137 -181 -12121 -147
rect -12053 -181 -12037 -147
rect -11979 -181 -11963 -147
rect -11895 -181 -11879 -147
rect -11821 -181 -11805 -147
rect -11737 -181 -11721 -147
rect -11663 -181 -11647 -147
rect -11579 -181 -11563 -147
rect -11505 -181 -11489 -147
rect -11421 -181 -11405 -147
rect -11347 -181 -11331 -147
rect -11263 -181 -11247 -147
rect -11189 -181 -11173 -147
rect -11105 -181 -11089 -147
rect -11031 -181 -11015 -147
rect -10947 -181 -10931 -147
rect -10873 -181 -10857 -147
rect -10789 -181 -10773 -147
rect -10715 -181 -10699 -147
rect -10631 -181 -10615 -147
rect -10557 -181 -10541 -147
rect -10473 -181 -10457 -147
rect -10399 -181 -10383 -147
rect -10315 -181 -10299 -147
rect -10241 -181 -10225 -147
rect -10157 -181 -10141 -147
rect -10083 -181 -10067 -147
rect -9999 -181 -9983 -147
rect -9925 -181 -9909 -147
rect -9841 -181 -9825 -147
rect -9767 -181 -9751 -147
rect -9683 -181 -9667 -147
rect -9609 -181 -9593 -147
rect -9525 -181 -9509 -147
rect -9451 -181 -9435 -147
rect -9367 -181 -9351 -147
rect -9293 -181 -9277 -147
rect -9209 -181 -9193 -147
rect -9135 -181 -9119 -147
rect -9051 -181 -9035 -147
rect -8977 -181 -8961 -147
rect -8893 -181 -8877 -147
rect -8819 -181 -8803 -147
rect -8735 -181 -8719 -147
rect -8661 -181 -8645 -147
rect -8577 -181 -8561 -147
rect -8503 -181 -8487 -147
rect -8419 -181 -8403 -147
rect -8345 -181 -8329 -147
rect -8261 -181 -8245 -147
rect -8187 -181 -8171 -147
rect -8103 -181 -8087 -147
rect -8029 -181 -8013 -147
rect -7945 -181 -7929 -147
rect -7871 -181 -7855 -147
rect -7787 -181 -7771 -147
rect -7713 -181 -7697 -147
rect -7629 -181 -7613 -147
rect -7555 -181 -7539 -147
rect -7471 -181 -7455 -147
rect -7397 -181 -7381 -147
rect -7313 -181 -7297 -147
rect -7239 -181 -7223 -147
rect -7155 -181 -7139 -147
rect -7081 -181 -7065 -147
rect -6997 -181 -6981 -147
rect -6923 -181 -6907 -147
rect -6839 -181 -6823 -147
rect -6765 -181 -6749 -147
rect -6681 -181 -6665 -147
rect -6607 -181 -6591 -147
rect -6523 -181 -6507 -147
rect -6449 -181 -6433 -147
rect -6365 -181 -6349 -147
rect -6291 -181 -6275 -147
rect -6207 -181 -6191 -147
rect -6133 -181 -6117 -147
rect -6049 -181 -6033 -147
rect -5975 -181 -5959 -147
rect -5891 -181 -5875 -147
rect -5817 -181 -5801 -147
rect -5733 -181 -5717 -147
rect -5659 -181 -5643 -147
rect -5575 -181 -5559 -147
rect -5501 -181 -5485 -147
rect -5417 -181 -5401 -147
rect -5343 -181 -5327 -147
rect -5259 -181 -5243 -147
rect -5185 -181 -5169 -147
rect -5101 -181 -5085 -147
rect -5027 -181 -5011 -147
rect -4943 -181 -4927 -147
rect -4869 -181 -4853 -147
rect -4785 -181 -4769 -147
rect -4711 -181 -4695 -147
rect -4627 -181 -4611 -147
rect -4553 -181 -4537 -147
rect -4469 -181 -4453 -147
rect -4395 -181 -4379 -147
rect -4311 -181 -4295 -147
rect -4237 -181 -4221 -147
rect -4153 -181 -4137 -147
rect -4079 -181 -4063 -147
rect -3995 -181 -3979 -147
rect -3921 -181 -3905 -147
rect -3837 -181 -3821 -147
rect -3763 -181 -3747 -147
rect -3679 -181 -3663 -147
rect -3605 -181 -3589 -147
rect -3521 -181 -3505 -147
rect -3447 -181 -3431 -147
rect -3363 -181 -3347 -147
rect -3289 -181 -3273 -147
rect -3205 -181 -3189 -147
rect -3131 -181 -3115 -147
rect -3047 -181 -3031 -147
rect -2973 -181 -2957 -147
rect -2889 -181 -2873 -147
rect -2815 -181 -2799 -147
rect -2731 -181 -2715 -147
rect -2657 -181 -2641 -147
rect -2573 -181 -2557 -147
rect -2499 -181 -2483 -147
rect -2415 -181 -2399 -147
rect -2341 -181 -2325 -147
rect -2257 -181 -2241 -147
rect -2183 -181 -2167 -147
rect -2099 -181 -2083 -147
rect -2025 -181 -2009 -147
rect -1941 -181 -1925 -147
rect -1867 -181 -1851 -147
rect -1783 -181 -1767 -147
rect -1709 -181 -1693 -147
rect -1625 -181 -1609 -147
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect 1609 -181 1625 -147
rect 1693 -181 1709 -147
rect 1767 -181 1783 -147
rect 1851 -181 1867 -147
rect 1925 -181 1941 -147
rect 2009 -181 2025 -147
rect 2083 -181 2099 -147
rect 2167 -181 2183 -147
rect 2241 -181 2257 -147
rect 2325 -181 2341 -147
rect 2399 -181 2415 -147
rect 2483 -181 2499 -147
rect 2557 -181 2573 -147
rect 2641 -181 2657 -147
rect 2715 -181 2731 -147
rect 2799 -181 2815 -147
rect 2873 -181 2889 -147
rect 2957 -181 2973 -147
rect 3031 -181 3047 -147
rect 3115 -181 3131 -147
rect 3189 -181 3205 -147
rect 3273 -181 3289 -147
rect 3347 -181 3363 -147
rect 3431 -181 3447 -147
rect 3505 -181 3521 -147
rect 3589 -181 3605 -147
rect 3663 -181 3679 -147
rect 3747 -181 3763 -147
rect 3821 -181 3837 -147
rect 3905 -181 3921 -147
rect 3979 -181 3995 -147
rect 4063 -181 4079 -147
rect 4137 -181 4153 -147
rect 4221 -181 4237 -147
rect 4295 -181 4311 -147
rect 4379 -181 4395 -147
rect 4453 -181 4469 -147
rect 4537 -181 4553 -147
rect 4611 -181 4627 -147
rect 4695 -181 4711 -147
rect 4769 -181 4785 -147
rect 4853 -181 4869 -147
rect 4927 -181 4943 -147
rect 5011 -181 5027 -147
rect 5085 -181 5101 -147
rect 5169 -181 5185 -147
rect 5243 -181 5259 -147
rect 5327 -181 5343 -147
rect 5401 -181 5417 -147
rect 5485 -181 5501 -147
rect 5559 -181 5575 -147
rect 5643 -181 5659 -147
rect 5717 -181 5733 -147
rect 5801 -181 5817 -147
rect 5875 -181 5891 -147
rect 5959 -181 5975 -147
rect 6033 -181 6049 -147
rect 6117 -181 6133 -147
rect 6191 -181 6207 -147
rect 6275 -181 6291 -147
rect 6349 -181 6365 -147
rect 6433 -181 6449 -147
rect 6507 -181 6523 -147
rect 6591 -181 6607 -147
rect 6665 -181 6681 -147
rect 6749 -181 6765 -147
rect 6823 -181 6839 -147
rect 6907 -181 6923 -147
rect 6981 -181 6997 -147
rect 7065 -181 7081 -147
rect 7139 -181 7155 -147
rect 7223 -181 7239 -147
rect 7297 -181 7313 -147
rect 7381 -181 7397 -147
rect 7455 -181 7471 -147
rect 7539 -181 7555 -147
rect 7613 -181 7629 -147
rect 7697 -181 7713 -147
rect 7771 -181 7787 -147
rect 7855 -181 7871 -147
rect 7929 -181 7945 -147
rect 8013 -181 8029 -147
rect 8087 -181 8103 -147
rect 8171 -181 8187 -147
rect 8245 -181 8261 -147
rect 8329 -181 8345 -147
rect 8403 -181 8419 -147
rect 8487 -181 8503 -147
rect 8561 -181 8577 -147
rect 8645 -181 8661 -147
rect 8719 -181 8735 -147
rect 8803 -181 8819 -147
rect 8877 -181 8893 -147
rect 8961 -181 8977 -147
rect 9035 -181 9051 -147
rect 9119 -181 9135 -147
rect 9193 -181 9209 -147
rect 9277 -181 9293 -147
rect 9351 -181 9367 -147
rect 9435 -181 9451 -147
rect 9509 -181 9525 -147
rect 9593 -181 9609 -147
rect 9667 -181 9683 -147
rect 9751 -181 9767 -147
rect 9825 -181 9841 -147
rect 9909 -181 9925 -147
rect 9983 -181 9999 -147
rect 10067 -181 10083 -147
rect 10141 -181 10157 -147
rect 10225 -181 10241 -147
rect 10299 -181 10315 -147
rect 10383 -181 10399 -147
rect 10457 -181 10473 -147
rect 10541 -181 10557 -147
rect 10615 -181 10631 -147
rect 10699 -181 10715 -147
rect 10773 -181 10789 -147
rect 10857 -181 10873 -147
rect 10931 -181 10947 -147
rect 11015 -181 11031 -147
rect 11089 -181 11105 -147
rect 11173 -181 11189 -147
rect 11247 -181 11263 -147
rect 11331 -181 11347 -147
rect 11405 -181 11421 -147
rect 11489 -181 11505 -147
rect 11563 -181 11579 -147
rect 11647 -181 11663 -147
rect 11721 -181 11737 -147
rect 11805 -181 11821 -147
rect 11879 -181 11895 -147
rect 11963 -181 11979 -147
rect 12037 -181 12053 -147
rect 12121 -181 12137 -147
rect 12195 -181 12211 -147
rect 12279 -181 12295 -147
rect 12353 -181 12369 -147
rect 12437 -181 12453 -147
rect 12511 -181 12527 -147
rect 12595 -181 12611 -147
rect 12669 -181 12685 -147
rect 12753 -181 12769 -147
rect 12827 -181 12843 -147
rect 12911 -181 12927 -147
rect 12985 -181 13001 -147
rect 13069 -181 13085 -147
rect 13143 -181 13159 -147
rect 13227 -181 13243 -147
rect 13301 -181 13317 -147
rect 13385 -181 13401 -147
rect 13459 -181 13475 -147
rect 13543 -181 13559 -147
rect 13617 -181 13633 -147
rect 13701 -181 13717 -147
rect 13775 -181 13791 -147
rect 13859 -181 13875 -147
rect 13933 -181 13949 -147
rect 14017 -181 14033 -147
rect 14091 -181 14107 -147
rect 14175 -181 14191 -147
rect 14249 -181 14265 -147
rect 14333 -181 14349 -147
rect 14407 -181 14423 -147
rect 14491 -181 14507 -147
rect 14565 -181 14581 -147
rect 14649 -181 14665 -147
rect 14723 -181 14739 -147
rect 14807 -181 14823 -147
rect 14881 -181 14897 -147
rect 14965 -181 14981 -147
rect 15039 -181 15055 -147
rect 15123 -181 15139 -147
rect 15197 -181 15213 -147
rect 15281 -181 15297 -147
rect 15355 -181 15371 -147
rect 15439 -181 15455 -147
rect 15513 -181 15529 -147
rect 15597 -181 15613 -147
rect 15671 -181 15687 -147
rect 15755 -181 15771 -147
rect -15951 -285 -15917 -223
rect 15917 -285 15951 -223
rect -15951 -319 -15855 -285
rect 15855 -319 15951 -285
<< viali >>
rect -15755 147 -15687 181
rect -15597 147 -15529 181
rect -15439 147 -15371 181
rect -15281 147 -15213 181
rect -15123 147 -15055 181
rect -14965 147 -14897 181
rect -14807 147 -14739 181
rect -14649 147 -14581 181
rect -14491 147 -14423 181
rect -14333 147 -14265 181
rect -14175 147 -14107 181
rect -14017 147 -13949 181
rect -13859 147 -13791 181
rect -13701 147 -13633 181
rect -13543 147 -13475 181
rect -13385 147 -13317 181
rect -13227 147 -13159 181
rect -13069 147 -13001 181
rect -12911 147 -12843 181
rect -12753 147 -12685 181
rect -12595 147 -12527 181
rect -12437 147 -12369 181
rect -12279 147 -12211 181
rect -12121 147 -12053 181
rect -11963 147 -11895 181
rect -11805 147 -11737 181
rect -11647 147 -11579 181
rect -11489 147 -11421 181
rect -11331 147 -11263 181
rect -11173 147 -11105 181
rect -11015 147 -10947 181
rect -10857 147 -10789 181
rect -10699 147 -10631 181
rect -10541 147 -10473 181
rect -10383 147 -10315 181
rect -10225 147 -10157 181
rect -10067 147 -9999 181
rect -9909 147 -9841 181
rect -9751 147 -9683 181
rect -9593 147 -9525 181
rect -9435 147 -9367 181
rect -9277 147 -9209 181
rect -9119 147 -9051 181
rect -8961 147 -8893 181
rect -8803 147 -8735 181
rect -8645 147 -8577 181
rect -8487 147 -8419 181
rect -8329 147 -8261 181
rect -8171 147 -8103 181
rect -8013 147 -7945 181
rect -7855 147 -7787 181
rect -7697 147 -7629 181
rect -7539 147 -7471 181
rect -7381 147 -7313 181
rect -7223 147 -7155 181
rect -7065 147 -6997 181
rect -6907 147 -6839 181
rect -6749 147 -6681 181
rect -6591 147 -6523 181
rect -6433 147 -6365 181
rect -6275 147 -6207 181
rect -6117 147 -6049 181
rect -5959 147 -5891 181
rect -5801 147 -5733 181
rect -5643 147 -5575 181
rect -5485 147 -5417 181
rect -5327 147 -5259 181
rect -5169 147 -5101 181
rect -5011 147 -4943 181
rect -4853 147 -4785 181
rect -4695 147 -4627 181
rect -4537 147 -4469 181
rect -4379 147 -4311 181
rect -4221 147 -4153 181
rect -4063 147 -3995 181
rect -3905 147 -3837 181
rect -3747 147 -3679 181
rect -3589 147 -3521 181
rect -3431 147 -3363 181
rect -3273 147 -3205 181
rect -3115 147 -3047 181
rect -2957 147 -2889 181
rect -2799 147 -2731 181
rect -2641 147 -2573 181
rect -2483 147 -2415 181
rect -2325 147 -2257 181
rect -2167 147 -2099 181
rect -2009 147 -1941 181
rect -1851 147 -1783 181
rect -1693 147 -1625 181
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect 1625 147 1693 181
rect 1783 147 1851 181
rect 1941 147 2009 181
rect 2099 147 2167 181
rect 2257 147 2325 181
rect 2415 147 2483 181
rect 2573 147 2641 181
rect 2731 147 2799 181
rect 2889 147 2957 181
rect 3047 147 3115 181
rect 3205 147 3273 181
rect 3363 147 3431 181
rect 3521 147 3589 181
rect 3679 147 3747 181
rect 3837 147 3905 181
rect 3995 147 4063 181
rect 4153 147 4221 181
rect 4311 147 4379 181
rect 4469 147 4537 181
rect 4627 147 4695 181
rect 4785 147 4853 181
rect 4943 147 5011 181
rect 5101 147 5169 181
rect 5259 147 5327 181
rect 5417 147 5485 181
rect 5575 147 5643 181
rect 5733 147 5801 181
rect 5891 147 5959 181
rect 6049 147 6117 181
rect 6207 147 6275 181
rect 6365 147 6433 181
rect 6523 147 6591 181
rect 6681 147 6749 181
rect 6839 147 6907 181
rect 6997 147 7065 181
rect 7155 147 7223 181
rect 7313 147 7381 181
rect 7471 147 7539 181
rect 7629 147 7697 181
rect 7787 147 7855 181
rect 7945 147 8013 181
rect 8103 147 8171 181
rect 8261 147 8329 181
rect 8419 147 8487 181
rect 8577 147 8645 181
rect 8735 147 8803 181
rect 8893 147 8961 181
rect 9051 147 9119 181
rect 9209 147 9277 181
rect 9367 147 9435 181
rect 9525 147 9593 181
rect 9683 147 9751 181
rect 9841 147 9909 181
rect 9999 147 10067 181
rect 10157 147 10225 181
rect 10315 147 10383 181
rect 10473 147 10541 181
rect 10631 147 10699 181
rect 10789 147 10857 181
rect 10947 147 11015 181
rect 11105 147 11173 181
rect 11263 147 11331 181
rect 11421 147 11489 181
rect 11579 147 11647 181
rect 11737 147 11805 181
rect 11895 147 11963 181
rect 12053 147 12121 181
rect 12211 147 12279 181
rect 12369 147 12437 181
rect 12527 147 12595 181
rect 12685 147 12753 181
rect 12843 147 12911 181
rect 13001 147 13069 181
rect 13159 147 13227 181
rect 13317 147 13385 181
rect 13475 147 13543 181
rect 13633 147 13701 181
rect 13791 147 13859 181
rect 13949 147 14017 181
rect 14107 147 14175 181
rect 14265 147 14333 181
rect 14423 147 14491 181
rect 14581 147 14649 181
rect 14739 147 14807 181
rect 14897 147 14965 181
rect 15055 147 15123 181
rect 15213 147 15281 181
rect 15371 147 15439 181
rect 15529 147 15597 181
rect 15687 147 15755 181
rect -15817 -88 -15783 88
rect -15659 -88 -15625 88
rect -15501 -88 -15467 88
rect -15343 -88 -15309 88
rect -15185 -88 -15151 88
rect -15027 -88 -14993 88
rect -14869 -88 -14835 88
rect -14711 -88 -14677 88
rect -14553 -88 -14519 88
rect -14395 -88 -14361 88
rect -14237 -88 -14203 88
rect -14079 -88 -14045 88
rect -13921 -88 -13887 88
rect -13763 -88 -13729 88
rect -13605 -88 -13571 88
rect -13447 -88 -13413 88
rect -13289 -88 -13255 88
rect -13131 -88 -13097 88
rect -12973 -88 -12939 88
rect -12815 -88 -12781 88
rect -12657 -88 -12623 88
rect -12499 -88 -12465 88
rect -12341 -88 -12307 88
rect -12183 -88 -12149 88
rect -12025 -88 -11991 88
rect -11867 -88 -11833 88
rect -11709 -88 -11675 88
rect -11551 -88 -11517 88
rect -11393 -88 -11359 88
rect -11235 -88 -11201 88
rect -11077 -88 -11043 88
rect -10919 -88 -10885 88
rect -10761 -88 -10727 88
rect -10603 -88 -10569 88
rect -10445 -88 -10411 88
rect -10287 -88 -10253 88
rect -10129 -88 -10095 88
rect -9971 -88 -9937 88
rect -9813 -88 -9779 88
rect -9655 -88 -9621 88
rect -9497 -88 -9463 88
rect -9339 -88 -9305 88
rect -9181 -88 -9147 88
rect -9023 -88 -8989 88
rect -8865 -88 -8831 88
rect -8707 -88 -8673 88
rect -8549 -88 -8515 88
rect -8391 -88 -8357 88
rect -8233 -88 -8199 88
rect -8075 -88 -8041 88
rect -7917 -88 -7883 88
rect -7759 -88 -7725 88
rect -7601 -88 -7567 88
rect -7443 -88 -7409 88
rect -7285 -88 -7251 88
rect -7127 -88 -7093 88
rect -6969 -88 -6935 88
rect -6811 -88 -6777 88
rect -6653 -88 -6619 88
rect -6495 -88 -6461 88
rect -6337 -88 -6303 88
rect -6179 -88 -6145 88
rect -6021 -88 -5987 88
rect -5863 -88 -5829 88
rect -5705 -88 -5671 88
rect -5547 -88 -5513 88
rect -5389 -88 -5355 88
rect -5231 -88 -5197 88
rect -5073 -88 -5039 88
rect -4915 -88 -4881 88
rect -4757 -88 -4723 88
rect -4599 -88 -4565 88
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect 4565 -88 4599 88
rect 4723 -88 4757 88
rect 4881 -88 4915 88
rect 5039 -88 5073 88
rect 5197 -88 5231 88
rect 5355 -88 5389 88
rect 5513 -88 5547 88
rect 5671 -88 5705 88
rect 5829 -88 5863 88
rect 5987 -88 6021 88
rect 6145 -88 6179 88
rect 6303 -88 6337 88
rect 6461 -88 6495 88
rect 6619 -88 6653 88
rect 6777 -88 6811 88
rect 6935 -88 6969 88
rect 7093 -88 7127 88
rect 7251 -88 7285 88
rect 7409 -88 7443 88
rect 7567 -88 7601 88
rect 7725 -88 7759 88
rect 7883 -88 7917 88
rect 8041 -88 8075 88
rect 8199 -88 8233 88
rect 8357 -88 8391 88
rect 8515 -88 8549 88
rect 8673 -88 8707 88
rect 8831 -88 8865 88
rect 8989 -88 9023 88
rect 9147 -88 9181 88
rect 9305 -88 9339 88
rect 9463 -88 9497 88
rect 9621 -88 9655 88
rect 9779 -88 9813 88
rect 9937 -88 9971 88
rect 10095 -88 10129 88
rect 10253 -88 10287 88
rect 10411 -88 10445 88
rect 10569 -88 10603 88
rect 10727 -88 10761 88
rect 10885 -88 10919 88
rect 11043 -88 11077 88
rect 11201 -88 11235 88
rect 11359 -88 11393 88
rect 11517 -88 11551 88
rect 11675 -88 11709 88
rect 11833 -88 11867 88
rect 11991 -88 12025 88
rect 12149 -88 12183 88
rect 12307 -88 12341 88
rect 12465 -88 12499 88
rect 12623 -88 12657 88
rect 12781 -88 12815 88
rect 12939 -88 12973 88
rect 13097 -88 13131 88
rect 13255 -88 13289 88
rect 13413 -88 13447 88
rect 13571 -88 13605 88
rect 13729 -88 13763 88
rect 13887 -88 13921 88
rect 14045 -88 14079 88
rect 14203 -88 14237 88
rect 14361 -88 14395 88
rect 14519 -88 14553 88
rect 14677 -88 14711 88
rect 14835 -88 14869 88
rect 14993 -88 15027 88
rect 15151 -88 15185 88
rect 15309 -88 15343 88
rect 15467 -88 15501 88
rect 15625 -88 15659 88
rect 15783 -88 15817 88
rect -15755 -181 -15687 -147
rect -15597 -181 -15529 -147
rect -15439 -181 -15371 -147
rect -15281 -181 -15213 -147
rect -15123 -181 -15055 -147
rect -14965 -181 -14897 -147
rect -14807 -181 -14739 -147
rect -14649 -181 -14581 -147
rect -14491 -181 -14423 -147
rect -14333 -181 -14265 -147
rect -14175 -181 -14107 -147
rect -14017 -181 -13949 -147
rect -13859 -181 -13791 -147
rect -13701 -181 -13633 -147
rect -13543 -181 -13475 -147
rect -13385 -181 -13317 -147
rect -13227 -181 -13159 -147
rect -13069 -181 -13001 -147
rect -12911 -181 -12843 -147
rect -12753 -181 -12685 -147
rect -12595 -181 -12527 -147
rect -12437 -181 -12369 -147
rect -12279 -181 -12211 -147
rect -12121 -181 -12053 -147
rect -11963 -181 -11895 -147
rect -11805 -181 -11737 -147
rect -11647 -181 -11579 -147
rect -11489 -181 -11421 -147
rect -11331 -181 -11263 -147
rect -11173 -181 -11105 -147
rect -11015 -181 -10947 -147
rect -10857 -181 -10789 -147
rect -10699 -181 -10631 -147
rect -10541 -181 -10473 -147
rect -10383 -181 -10315 -147
rect -10225 -181 -10157 -147
rect -10067 -181 -9999 -147
rect -9909 -181 -9841 -147
rect -9751 -181 -9683 -147
rect -9593 -181 -9525 -147
rect -9435 -181 -9367 -147
rect -9277 -181 -9209 -147
rect -9119 -181 -9051 -147
rect -8961 -181 -8893 -147
rect -8803 -181 -8735 -147
rect -8645 -181 -8577 -147
rect -8487 -181 -8419 -147
rect -8329 -181 -8261 -147
rect -8171 -181 -8103 -147
rect -8013 -181 -7945 -147
rect -7855 -181 -7787 -147
rect -7697 -181 -7629 -147
rect -7539 -181 -7471 -147
rect -7381 -181 -7313 -147
rect -7223 -181 -7155 -147
rect -7065 -181 -6997 -147
rect -6907 -181 -6839 -147
rect -6749 -181 -6681 -147
rect -6591 -181 -6523 -147
rect -6433 -181 -6365 -147
rect -6275 -181 -6207 -147
rect -6117 -181 -6049 -147
rect -5959 -181 -5891 -147
rect -5801 -181 -5733 -147
rect -5643 -181 -5575 -147
rect -5485 -181 -5417 -147
rect -5327 -181 -5259 -147
rect -5169 -181 -5101 -147
rect -5011 -181 -4943 -147
rect -4853 -181 -4785 -147
rect -4695 -181 -4627 -147
rect -4537 -181 -4469 -147
rect -4379 -181 -4311 -147
rect -4221 -181 -4153 -147
rect -4063 -181 -3995 -147
rect -3905 -181 -3837 -147
rect -3747 -181 -3679 -147
rect -3589 -181 -3521 -147
rect -3431 -181 -3363 -147
rect -3273 -181 -3205 -147
rect -3115 -181 -3047 -147
rect -2957 -181 -2889 -147
rect -2799 -181 -2731 -147
rect -2641 -181 -2573 -147
rect -2483 -181 -2415 -147
rect -2325 -181 -2257 -147
rect -2167 -181 -2099 -147
rect -2009 -181 -1941 -147
rect -1851 -181 -1783 -147
rect -1693 -181 -1625 -147
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
rect 1625 -181 1693 -147
rect 1783 -181 1851 -147
rect 1941 -181 2009 -147
rect 2099 -181 2167 -147
rect 2257 -181 2325 -147
rect 2415 -181 2483 -147
rect 2573 -181 2641 -147
rect 2731 -181 2799 -147
rect 2889 -181 2957 -147
rect 3047 -181 3115 -147
rect 3205 -181 3273 -147
rect 3363 -181 3431 -147
rect 3521 -181 3589 -147
rect 3679 -181 3747 -147
rect 3837 -181 3905 -147
rect 3995 -181 4063 -147
rect 4153 -181 4221 -147
rect 4311 -181 4379 -147
rect 4469 -181 4537 -147
rect 4627 -181 4695 -147
rect 4785 -181 4853 -147
rect 4943 -181 5011 -147
rect 5101 -181 5169 -147
rect 5259 -181 5327 -147
rect 5417 -181 5485 -147
rect 5575 -181 5643 -147
rect 5733 -181 5801 -147
rect 5891 -181 5959 -147
rect 6049 -181 6117 -147
rect 6207 -181 6275 -147
rect 6365 -181 6433 -147
rect 6523 -181 6591 -147
rect 6681 -181 6749 -147
rect 6839 -181 6907 -147
rect 6997 -181 7065 -147
rect 7155 -181 7223 -147
rect 7313 -181 7381 -147
rect 7471 -181 7539 -147
rect 7629 -181 7697 -147
rect 7787 -181 7855 -147
rect 7945 -181 8013 -147
rect 8103 -181 8171 -147
rect 8261 -181 8329 -147
rect 8419 -181 8487 -147
rect 8577 -181 8645 -147
rect 8735 -181 8803 -147
rect 8893 -181 8961 -147
rect 9051 -181 9119 -147
rect 9209 -181 9277 -147
rect 9367 -181 9435 -147
rect 9525 -181 9593 -147
rect 9683 -181 9751 -147
rect 9841 -181 9909 -147
rect 9999 -181 10067 -147
rect 10157 -181 10225 -147
rect 10315 -181 10383 -147
rect 10473 -181 10541 -147
rect 10631 -181 10699 -147
rect 10789 -181 10857 -147
rect 10947 -181 11015 -147
rect 11105 -181 11173 -147
rect 11263 -181 11331 -147
rect 11421 -181 11489 -147
rect 11579 -181 11647 -147
rect 11737 -181 11805 -147
rect 11895 -181 11963 -147
rect 12053 -181 12121 -147
rect 12211 -181 12279 -147
rect 12369 -181 12437 -147
rect 12527 -181 12595 -147
rect 12685 -181 12753 -147
rect 12843 -181 12911 -147
rect 13001 -181 13069 -147
rect 13159 -181 13227 -147
rect 13317 -181 13385 -147
rect 13475 -181 13543 -147
rect 13633 -181 13701 -147
rect 13791 -181 13859 -147
rect 13949 -181 14017 -147
rect 14107 -181 14175 -147
rect 14265 -181 14333 -147
rect 14423 -181 14491 -147
rect 14581 -181 14649 -147
rect 14739 -181 14807 -147
rect 14897 -181 14965 -147
rect 15055 -181 15123 -147
rect 15213 -181 15281 -147
rect 15371 -181 15439 -147
rect 15529 -181 15597 -147
rect 15687 -181 15755 -147
<< metal1 >>
rect -15767 181 -15675 187
rect -15767 147 -15755 181
rect -15687 147 -15675 181
rect -15767 141 -15675 147
rect -15609 181 -15517 187
rect -15609 147 -15597 181
rect -15529 147 -15517 181
rect -15609 141 -15517 147
rect -15451 181 -15359 187
rect -15451 147 -15439 181
rect -15371 147 -15359 181
rect -15451 141 -15359 147
rect -15293 181 -15201 187
rect -15293 147 -15281 181
rect -15213 147 -15201 181
rect -15293 141 -15201 147
rect -15135 181 -15043 187
rect -15135 147 -15123 181
rect -15055 147 -15043 181
rect -15135 141 -15043 147
rect -14977 181 -14885 187
rect -14977 147 -14965 181
rect -14897 147 -14885 181
rect -14977 141 -14885 147
rect -14819 181 -14727 187
rect -14819 147 -14807 181
rect -14739 147 -14727 181
rect -14819 141 -14727 147
rect -14661 181 -14569 187
rect -14661 147 -14649 181
rect -14581 147 -14569 181
rect -14661 141 -14569 147
rect -14503 181 -14411 187
rect -14503 147 -14491 181
rect -14423 147 -14411 181
rect -14503 141 -14411 147
rect -14345 181 -14253 187
rect -14345 147 -14333 181
rect -14265 147 -14253 181
rect -14345 141 -14253 147
rect -14187 181 -14095 187
rect -14187 147 -14175 181
rect -14107 147 -14095 181
rect -14187 141 -14095 147
rect -14029 181 -13937 187
rect -14029 147 -14017 181
rect -13949 147 -13937 181
rect -14029 141 -13937 147
rect -13871 181 -13779 187
rect -13871 147 -13859 181
rect -13791 147 -13779 181
rect -13871 141 -13779 147
rect -13713 181 -13621 187
rect -13713 147 -13701 181
rect -13633 147 -13621 181
rect -13713 141 -13621 147
rect -13555 181 -13463 187
rect -13555 147 -13543 181
rect -13475 147 -13463 181
rect -13555 141 -13463 147
rect -13397 181 -13305 187
rect -13397 147 -13385 181
rect -13317 147 -13305 181
rect -13397 141 -13305 147
rect -13239 181 -13147 187
rect -13239 147 -13227 181
rect -13159 147 -13147 181
rect -13239 141 -13147 147
rect -13081 181 -12989 187
rect -13081 147 -13069 181
rect -13001 147 -12989 181
rect -13081 141 -12989 147
rect -12923 181 -12831 187
rect -12923 147 -12911 181
rect -12843 147 -12831 181
rect -12923 141 -12831 147
rect -12765 181 -12673 187
rect -12765 147 -12753 181
rect -12685 147 -12673 181
rect -12765 141 -12673 147
rect -12607 181 -12515 187
rect -12607 147 -12595 181
rect -12527 147 -12515 181
rect -12607 141 -12515 147
rect -12449 181 -12357 187
rect -12449 147 -12437 181
rect -12369 147 -12357 181
rect -12449 141 -12357 147
rect -12291 181 -12199 187
rect -12291 147 -12279 181
rect -12211 147 -12199 181
rect -12291 141 -12199 147
rect -12133 181 -12041 187
rect -12133 147 -12121 181
rect -12053 147 -12041 181
rect -12133 141 -12041 147
rect -11975 181 -11883 187
rect -11975 147 -11963 181
rect -11895 147 -11883 181
rect -11975 141 -11883 147
rect -11817 181 -11725 187
rect -11817 147 -11805 181
rect -11737 147 -11725 181
rect -11817 141 -11725 147
rect -11659 181 -11567 187
rect -11659 147 -11647 181
rect -11579 147 -11567 181
rect -11659 141 -11567 147
rect -11501 181 -11409 187
rect -11501 147 -11489 181
rect -11421 147 -11409 181
rect -11501 141 -11409 147
rect -11343 181 -11251 187
rect -11343 147 -11331 181
rect -11263 147 -11251 181
rect -11343 141 -11251 147
rect -11185 181 -11093 187
rect -11185 147 -11173 181
rect -11105 147 -11093 181
rect -11185 141 -11093 147
rect -11027 181 -10935 187
rect -11027 147 -11015 181
rect -10947 147 -10935 181
rect -11027 141 -10935 147
rect -10869 181 -10777 187
rect -10869 147 -10857 181
rect -10789 147 -10777 181
rect -10869 141 -10777 147
rect -10711 181 -10619 187
rect -10711 147 -10699 181
rect -10631 147 -10619 181
rect -10711 141 -10619 147
rect -10553 181 -10461 187
rect -10553 147 -10541 181
rect -10473 147 -10461 181
rect -10553 141 -10461 147
rect -10395 181 -10303 187
rect -10395 147 -10383 181
rect -10315 147 -10303 181
rect -10395 141 -10303 147
rect -10237 181 -10145 187
rect -10237 147 -10225 181
rect -10157 147 -10145 181
rect -10237 141 -10145 147
rect -10079 181 -9987 187
rect -10079 147 -10067 181
rect -9999 147 -9987 181
rect -10079 141 -9987 147
rect -9921 181 -9829 187
rect -9921 147 -9909 181
rect -9841 147 -9829 181
rect -9921 141 -9829 147
rect -9763 181 -9671 187
rect -9763 147 -9751 181
rect -9683 147 -9671 181
rect -9763 141 -9671 147
rect -9605 181 -9513 187
rect -9605 147 -9593 181
rect -9525 147 -9513 181
rect -9605 141 -9513 147
rect -9447 181 -9355 187
rect -9447 147 -9435 181
rect -9367 147 -9355 181
rect -9447 141 -9355 147
rect -9289 181 -9197 187
rect -9289 147 -9277 181
rect -9209 147 -9197 181
rect -9289 141 -9197 147
rect -9131 181 -9039 187
rect -9131 147 -9119 181
rect -9051 147 -9039 181
rect -9131 141 -9039 147
rect -8973 181 -8881 187
rect -8973 147 -8961 181
rect -8893 147 -8881 181
rect -8973 141 -8881 147
rect -8815 181 -8723 187
rect -8815 147 -8803 181
rect -8735 147 -8723 181
rect -8815 141 -8723 147
rect -8657 181 -8565 187
rect -8657 147 -8645 181
rect -8577 147 -8565 181
rect -8657 141 -8565 147
rect -8499 181 -8407 187
rect -8499 147 -8487 181
rect -8419 147 -8407 181
rect -8499 141 -8407 147
rect -8341 181 -8249 187
rect -8341 147 -8329 181
rect -8261 147 -8249 181
rect -8341 141 -8249 147
rect -8183 181 -8091 187
rect -8183 147 -8171 181
rect -8103 147 -8091 181
rect -8183 141 -8091 147
rect -8025 181 -7933 187
rect -8025 147 -8013 181
rect -7945 147 -7933 181
rect -8025 141 -7933 147
rect -7867 181 -7775 187
rect -7867 147 -7855 181
rect -7787 147 -7775 181
rect -7867 141 -7775 147
rect -7709 181 -7617 187
rect -7709 147 -7697 181
rect -7629 147 -7617 181
rect -7709 141 -7617 147
rect -7551 181 -7459 187
rect -7551 147 -7539 181
rect -7471 147 -7459 181
rect -7551 141 -7459 147
rect -7393 181 -7301 187
rect -7393 147 -7381 181
rect -7313 147 -7301 181
rect -7393 141 -7301 147
rect -7235 181 -7143 187
rect -7235 147 -7223 181
rect -7155 147 -7143 181
rect -7235 141 -7143 147
rect -7077 181 -6985 187
rect -7077 147 -7065 181
rect -6997 147 -6985 181
rect -7077 141 -6985 147
rect -6919 181 -6827 187
rect -6919 147 -6907 181
rect -6839 147 -6827 181
rect -6919 141 -6827 147
rect -6761 181 -6669 187
rect -6761 147 -6749 181
rect -6681 147 -6669 181
rect -6761 141 -6669 147
rect -6603 181 -6511 187
rect -6603 147 -6591 181
rect -6523 147 -6511 181
rect -6603 141 -6511 147
rect -6445 181 -6353 187
rect -6445 147 -6433 181
rect -6365 147 -6353 181
rect -6445 141 -6353 147
rect -6287 181 -6195 187
rect -6287 147 -6275 181
rect -6207 147 -6195 181
rect -6287 141 -6195 147
rect -6129 181 -6037 187
rect -6129 147 -6117 181
rect -6049 147 -6037 181
rect -6129 141 -6037 147
rect -5971 181 -5879 187
rect -5971 147 -5959 181
rect -5891 147 -5879 181
rect -5971 141 -5879 147
rect -5813 181 -5721 187
rect -5813 147 -5801 181
rect -5733 147 -5721 181
rect -5813 141 -5721 147
rect -5655 181 -5563 187
rect -5655 147 -5643 181
rect -5575 147 -5563 181
rect -5655 141 -5563 147
rect -5497 181 -5405 187
rect -5497 147 -5485 181
rect -5417 147 -5405 181
rect -5497 141 -5405 147
rect -5339 181 -5247 187
rect -5339 147 -5327 181
rect -5259 147 -5247 181
rect -5339 141 -5247 147
rect -5181 181 -5089 187
rect -5181 147 -5169 181
rect -5101 147 -5089 181
rect -5181 141 -5089 147
rect -5023 181 -4931 187
rect -5023 147 -5011 181
rect -4943 147 -4931 181
rect -5023 141 -4931 147
rect -4865 181 -4773 187
rect -4865 147 -4853 181
rect -4785 147 -4773 181
rect -4865 141 -4773 147
rect -4707 181 -4615 187
rect -4707 147 -4695 181
rect -4627 147 -4615 181
rect -4707 141 -4615 147
rect -4549 181 -4457 187
rect -4549 147 -4537 181
rect -4469 147 -4457 181
rect -4549 141 -4457 147
rect -4391 181 -4299 187
rect -4391 147 -4379 181
rect -4311 147 -4299 181
rect -4391 141 -4299 147
rect -4233 181 -4141 187
rect -4233 147 -4221 181
rect -4153 147 -4141 181
rect -4233 141 -4141 147
rect -4075 181 -3983 187
rect -4075 147 -4063 181
rect -3995 147 -3983 181
rect -4075 141 -3983 147
rect -3917 181 -3825 187
rect -3917 147 -3905 181
rect -3837 147 -3825 181
rect -3917 141 -3825 147
rect -3759 181 -3667 187
rect -3759 147 -3747 181
rect -3679 147 -3667 181
rect -3759 141 -3667 147
rect -3601 181 -3509 187
rect -3601 147 -3589 181
rect -3521 147 -3509 181
rect -3601 141 -3509 147
rect -3443 181 -3351 187
rect -3443 147 -3431 181
rect -3363 147 -3351 181
rect -3443 141 -3351 147
rect -3285 181 -3193 187
rect -3285 147 -3273 181
rect -3205 147 -3193 181
rect -3285 141 -3193 147
rect -3127 181 -3035 187
rect -3127 147 -3115 181
rect -3047 147 -3035 181
rect -3127 141 -3035 147
rect -2969 181 -2877 187
rect -2969 147 -2957 181
rect -2889 147 -2877 181
rect -2969 141 -2877 147
rect -2811 181 -2719 187
rect -2811 147 -2799 181
rect -2731 147 -2719 181
rect -2811 141 -2719 147
rect -2653 181 -2561 187
rect -2653 147 -2641 181
rect -2573 147 -2561 181
rect -2653 141 -2561 147
rect -2495 181 -2403 187
rect -2495 147 -2483 181
rect -2415 147 -2403 181
rect -2495 141 -2403 147
rect -2337 181 -2245 187
rect -2337 147 -2325 181
rect -2257 147 -2245 181
rect -2337 141 -2245 147
rect -2179 181 -2087 187
rect -2179 147 -2167 181
rect -2099 147 -2087 181
rect -2179 141 -2087 147
rect -2021 181 -1929 187
rect -2021 147 -2009 181
rect -1941 147 -1929 181
rect -2021 141 -1929 147
rect -1863 181 -1771 187
rect -1863 147 -1851 181
rect -1783 147 -1771 181
rect -1863 141 -1771 147
rect -1705 181 -1613 187
rect -1705 147 -1693 181
rect -1625 147 -1613 181
rect -1705 141 -1613 147
rect -1547 181 -1455 187
rect -1547 147 -1535 181
rect -1467 147 -1455 181
rect -1547 141 -1455 147
rect -1389 181 -1297 187
rect -1389 147 -1377 181
rect -1309 147 -1297 181
rect -1389 141 -1297 147
rect -1231 181 -1139 187
rect -1231 147 -1219 181
rect -1151 147 -1139 181
rect -1231 141 -1139 147
rect -1073 181 -981 187
rect -1073 147 -1061 181
rect -993 147 -981 181
rect -1073 141 -981 147
rect -915 181 -823 187
rect -915 147 -903 181
rect -835 147 -823 181
rect -915 141 -823 147
rect -757 181 -665 187
rect -757 147 -745 181
rect -677 147 -665 181
rect -757 141 -665 147
rect -599 181 -507 187
rect -599 147 -587 181
rect -519 147 -507 181
rect -599 141 -507 147
rect -441 181 -349 187
rect -441 147 -429 181
rect -361 147 -349 181
rect -441 141 -349 147
rect -283 181 -191 187
rect -283 147 -271 181
rect -203 147 -191 181
rect -283 141 -191 147
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect 191 181 283 187
rect 191 147 203 181
rect 271 147 283 181
rect 191 141 283 147
rect 349 181 441 187
rect 349 147 361 181
rect 429 147 441 181
rect 349 141 441 147
rect 507 181 599 187
rect 507 147 519 181
rect 587 147 599 181
rect 507 141 599 147
rect 665 181 757 187
rect 665 147 677 181
rect 745 147 757 181
rect 665 141 757 147
rect 823 181 915 187
rect 823 147 835 181
rect 903 147 915 181
rect 823 141 915 147
rect 981 181 1073 187
rect 981 147 993 181
rect 1061 147 1073 181
rect 981 141 1073 147
rect 1139 181 1231 187
rect 1139 147 1151 181
rect 1219 147 1231 181
rect 1139 141 1231 147
rect 1297 181 1389 187
rect 1297 147 1309 181
rect 1377 147 1389 181
rect 1297 141 1389 147
rect 1455 181 1547 187
rect 1455 147 1467 181
rect 1535 147 1547 181
rect 1455 141 1547 147
rect 1613 181 1705 187
rect 1613 147 1625 181
rect 1693 147 1705 181
rect 1613 141 1705 147
rect 1771 181 1863 187
rect 1771 147 1783 181
rect 1851 147 1863 181
rect 1771 141 1863 147
rect 1929 181 2021 187
rect 1929 147 1941 181
rect 2009 147 2021 181
rect 1929 141 2021 147
rect 2087 181 2179 187
rect 2087 147 2099 181
rect 2167 147 2179 181
rect 2087 141 2179 147
rect 2245 181 2337 187
rect 2245 147 2257 181
rect 2325 147 2337 181
rect 2245 141 2337 147
rect 2403 181 2495 187
rect 2403 147 2415 181
rect 2483 147 2495 181
rect 2403 141 2495 147
rect 2561 181 2653 187
rect 2561 147 2573 181
rect 2641 147 2653 181
rect 2561 141 2653 147
rect 2719 181 2811 187
rect 2719 147 2731 181
rect 2799 147 2811 181
rect 2719 141 2811 147
rect 2877 181 2969 187
rect 2877 147 2889 181
rect 2957 147 2969 181
rect 2877 141 2969 147
rect 3035 181 3127 187
rect 3035 147 3047 181
rect 3115 147 3127 181
rect 3035 141 3127 147
rect 3193 181 3285 187
rect 3193 147 3205 181
rect 3273 147 3285 181
rect 3193 141 3285 147
rect 3351 181 3443 187
rect 3351 147 3363 181
rect 3431 147 3443 181
rect 3351 141 3443 147
rect 3509 181 3601 187
rect 3509 147 3521 181
rect 3589 147 3601 181
rect 3509 141 3601 147
rect 3667 181 3759 187
rect 3667 147 3679 181
rect 3747 147 3759 181
rect 3667 141 3759 147
rect 3825 181 3917 187
rect 3825 147 3837 181
rect 3905 147 3917 181
rect 3825 141 3917 147
rect 3983 181 4075 187
rect 3983 147 3995 181
rect 4063 147 4075 181
rect 3983 141 4075 147
rect 4141 181 4233 187
rect 4141 147 4153 181
rect 4221 147 4233 181
rect 4141 141 4233 147
rect 4299 181 4391 187
rect 4299 147 4311 181
rect 4379 147 4391 181
rect 4299 141 4391 147
rect 4457 181 4549 187
rect 4457 147 4469 181
rect 4537 147 4549 181
rect 4457 141 4549 147
rect 4615 181 4707 187
rect 4615 147 4627 181
rect 4695 147 4707 181
rect 4615 141 4707 147
rect 4773 181 4865 187
rect 4773 147 4785 181
rect 4853 147 4865 181
rect 4773 141 4865 147
rect 4931 181 5023 187
rect 4931 147 4943 181
rect 5011 147 5023 181
rect 4931 141 5023 147
rect 5089 181 5181 187
rect 5089 147 5101 181
rect 5169 147 5181 181
rect 5089 141 5181 147
rect 5247 181 5339 187
rect 5247 147 5259 181
rect 5327 147 5339 181
rect 5247 141 5339 147
rect 5405 181 5497 187
rect 5405 147 5417 181
rect 5485 147 5497 181
rect 5405 141 5497 147
rect 5563 181 5655 187
rect 5563 147 5575 181
rect 5643 147 5655 181
rect 5563 141 5655 147
rect 5721 181 5813 187
rect 5721 147 5733 181
rect 5801 147 5813 181
rect 5721 141 5813 147
rect 5879 181 5971 187
rect 5879 147 5891 181
rect 5959 147 5971 181
rect 5879 141 5971 147
rect 6037 181 6129 187
rect 6037 147 6049 181
rect 6117 147 6129 181
rect 6037 141 6129 147
rect 6195 181 6287 187
rect 6195 147 6207 181
rect 6275 147 6287 181
rect 6195 141 6287 147
rect 6353 181 6445 187
rect 6353 147 6365 181
rect 6433 147 6445 181
rect 6353 141 6445 147
rect 6511 181 6603 187
rect 6511 147 6523 181
rect 6591 147 6603 181
rect 6511 141 6603 147
rect 6669 181 6761 187
rect 6669 147 6681 181
rect 6749 147 6761 181
rect 6669 141 6761 147
rect 6827 181 6919 187
rect 6827 147 6839 181
rect 6907 147 6919 181
rect 6827 141 6919 147
rect 6985 181 7077 187
rect 6985 147 6997 181
rect 7065 147 7077 181
rect 6985 141 7077 147
rect 7143 181 7235 187
rect 7143 147 7155 181
rect 7223 147 7235 181
rect 7143 141 7235 147
rect 7301 181 7393 187
rect 7301 147 7313 181
rect 7381 147 7393 181
rect 7301 141 7393 147
rect 7459 181 7551 187
rect 7459 147 7471 181
rect 7539 147 7551 181
rect 7459 141 7551 147
rect 7617 181 7709 187
rect 7617 147 7629 181
rect 7697 147 7709 181
rect 7617 141 7709 147
rect 7775 181 7867 187
rect 7775 147 7787 181
rect 7855 147 7867 181
rect 7775 141 7867 147
rect 7933 181 8025 187
rect 7933 147 7945 181
rect 8013 147 8025 181
rect 7933 141 8025 147
rect 8091 181 8183 187
rect 8091 147 8103 181
rect 8171 147 8183 181
rect 8091 141 8183 147
rect 8249 181 8341 187
rect 8249 147 8261 181
rect 8329 147 8341 181
rect 8249 141 8341 147
rect 8407 181 8499 187
rect 8407 147 8419 181
rect 8487 147 8499 181
rect 8407 141 8499 147
rect 8565 181 8657 187
rect 8565 147 8577 181
rect 8645 147 8657 181
rect 8565 141 8657 147
rect 8723 181 8815 187
rect 8723 147 8735 181
rect 8803 147 8815 181
rect 8723 141 8815 147
rect 8881 181 8973 187
rect 8881 147 8893 181
rect 8961 147 8973 181
rect 8881 141 8973 147
rect 9039 181 9131 187
rect 9039 147 9051 181
rect 9119 147 9131 181
rect 9039 141 9131 147
rect 9197 181 9289 187
rect 9197 147 9209 181
rect 9277 147 9289 181
rect 9197 141 9289 147
rect 9355 181 9447 187
rect 9355 147 9367 181
rect 9435 147 9447 181
rect 9355 141 9447 147
rect 9513 181 9605 187
rect 9513 147 9525 181
rect 9593 147 9605 181
rect 9513 141 9605 147
rect 9671 181 9763 187
rect 9671 147 9683 181
rect 9751 147 9763 181
rect 9671 141 9763 147
rect 9829 181 9921 187
rect 9829 147 9841 181
rect 9909 147 9921 181
rect 9829 141 9921 147
rect 9987 181 10079 187
rect 9987 147 9999 181
rect 10067 147 10079 181
rect 9987 141 10079 147
rect 10145 181 10237 187
rect 10145 147 10157 181
rect 10225 147 10237 181
rect 10145 141 10237 147
rect 10303 181 10395 187
rect 10303 147 10315 181
rect 10383 147 10395 181
rect 10303 141 10395 147
rect 10461 181 10553 187
rect 10461 147 10473 181
rect 10541 147 10553 181
rect 10461 141 10553 147
rect 10619 181 10711 187
rect 10619 147 10631 181
rect 10699 147 10711 181
rect 10619 141 10711 147
rect 10777 181 10869 187
rect 10777 147 10789 181
rect 10857 147 10869 181
rect 10777 141 10869 147
rect 10935 181 11027 187
rect 10935 147 10947 181
rect 11015 147 11027 181
rect 10935 141 11027 147
rect 11093 181 11185 187
rect 11093 147 11105 181
rect 11173 147 11185 181
rect 11093 141 11185 147
rect 11251 181 11343 187
rect 11251 147 11263 181
rect 11331 147 11343 181
rect 11251 141 11343 147
rect 11409 181 11501 187
rect 11409 147 11421 181
rect 11489 147 11501 181
rect 11409 141 11501 147
rect 11567 181 11659 187
rect 11567 147 11579 181
rect 11647 147 11659 181
rect 11567 141 11659 147
rect 11725 181 11817 187
rect 11725 147 11737 181
rect 11805 147 11817 181
rect 11725 141 11817 147
rect 11883 181 11975 187
rect 11883 147 11895 181
rect 11963 147 11975 181
rect 11883 141 11975 147
rect 12041 181 12133 187
rect 12041 147 12053 181
rect 12121 147 12133 181
rect 12041 141 12133 147
rect 12199 181 12291 187
rect 12199 147 12211 181
rect 12279 147 12291 181
rect 12199 141 12291 147
rect 12357 181 12449 187
rect 12357 147 12369 181
rect 12437 147 12449 181
rect 12357 141 12449 147
rect 12515 181 12607 187
rect 12515 147 12527 181
rect 12595 147 12607 181
rect 12515 141 12607 147
rect 12673 181 12765 187
rect 12673 147 12685 181
rect 12753 147 12765 181
rect 12673 141 12765 147
rect 12831 181 12923 187
rect 12831 147 12843 181
rect 12911 147 12923 181
rect 12831 141 12923 147
rect 12989 181 13081 187
rect 12989 147 13001 181
rect 13069 147 13081 181
rect 12989 141 13081 147
rect 13147 181 13239 187
rect 13147 147 13159 181
rect 13227 147 13239 181
rect 13147 141 13239 147
rect 13305 181 13397 187
rect 13305 147 13317 181
rect 13385 147 13397 181
rect 13305 141 13397 147
rect 13463 181 13555 187
rect 13463 147 13475 181
rect 13543 147 13555 181
rect 13463 141 13555 147
rect 13621 181 13713 187
rect 13621 147 13633 181
rect 13701 147 13713 181
rect 13621 141 13713 147
rect 13779 181 13871 187
rect 13779 147 13791 181
rect 13859 147 13871 181
rect 13779 141 13871 147
rect 13937 181 14029 187
rect 13937 147 13949 181
rect 14017 147 14029 181
rect 13937 141 14029 147
rect 14095 181 14187 187
rect 14095 147 14107 181
rect 14175 147 14187 181
rect 14095 141 14187 147
rect 14253 181 14345 187
rect 14253 147 14265 181
rect 14333 147 14345 181
rect 14253 141 14345 147
rect 14411 181 14503 187
rect 14411 147 14423 181
rect 14491 147 14503 181
rect 14411 141 14503 147
rect 14569 181 14661 187
rect 14569 147 14581 181
rect 14649 147 14661 181
rect 14569 141 14661 147
rect 14727 181 14819 187
rect 14727 147 14739 181
rect 14807 147 14819 181
rect 14727 141 14819 147
rect 14885 181 14977 187
rect 14885 147 14897 181
rect 14965 147 14977 181
rect 14885 141 14977 147
rect 15043 181 15135 187
rect 15043 147 15055 181
rect 15123 147 15135 181
rect 15043 141 15135 147
rect 15201 181 15293 187
rect 15201 147 15213 181
rect 15281 147 15293 181
rect 15201 141 15293 147
rect 15359 181 15451 187
rect 15359 147 15371 181
rect 15439 147 15451 181
rect 15359 141 15451 147
rect 15517 181 15609 187
rect 15517 147 15529 181
rect 15597 147 15609 181
rect 15517 141 15609 147
rect 15675 181 15767 187
rect 15675 147 15687 181
rect 15755 147 15767 181
rect 15675 141 15767 147
rect -15823 88 -15777 100
rect -15823 -88 -15817 88
rect -15783 -88 -15777 88
rect -15823 -100 -15777 -88
rect -15665 88 -15619 100
rect -15665 -88 -15659 88
rect -15625 -88 -15619 88
rect -15665 -100 -15619 -88
rect -15507 88 -15461 100
rect -15507 -88 -15501 88
rect -15467 -88 -15461 88
rect -15507 -100 -15461 -88
rect -15349 88 -15303 100
rect -15349 -88 -15343 88
rect -15309 -88 -15303 88
rect -15349 -100 -15303 -88
rect -15191 88 -15145 100
rect -15191 -88 -15185 88
rect -15151 -88 -15145 88
rect -15191 -100 -15145 -88
rect -15033 88 -14987 100
rect -15033 -88 -15027 88
rect -14993 -88 -14987 88
rect -15033 -100 -14987 -88
rect -14875 88 -14829 100
rect -14875 -88 -14869 88
rect -14835 -88 -14829 88
rect -14875 -100 -14829 -88
rect -14717 88 -14671 100
rect -14717 -88 -14711 88
rect -14677 -88 -14671 88
rect -14717 -100 -14671 -88
rect -14559 88 -14513 100
rect -14559 -88 -14553 88
rect -14519 -88 -14513 88
rect -14559 -100 -14513 -88
rect -14401 88 -14355 100
rect -14401 -88 -14395 88
rect -14361 -88 -14355 88
rect -14401 -100 -14355 -88
rect -14243 88 -14197 100
rect -14243 -88 -14237 88
rect -14203 -88 -14197 88
rect -14243 -100 -14197 -88
rect -14085 88 -14039 100
rect -14085 -88 -14079 88
rect -14045 -88 -14039 88
rect -14085 -100 -14039 -88
rect -13927 88 -13881 100
rect -13927 -88 -13921 88
rect -13887 -88 -13881 88
rect -13927 -100 -13881 -88
rect -13769 88 -13723 100
rect -13769 -88 -13763 88
rect -13729 -88 -13723 88
rect -13769 -100 -13723 -88
rect -13611 88 -13565 100
rect -13611 -88 -13605 88
rect -13571 -88 -13565 88
rect -13611 -100 -13565 -88
rect -13453 88 -13407 100
rect -13453 -88 -13447 88
rect -13413 -88 -13407 88
rect -13453 -100 -13407 -88
rect -13295 88 -13249 100
rect -13295 -88 -13289 88
rect -13255 -88 -13249 88
rect -13295 -100 -13249 -88
rect -13137 88 -13091 100
rect -13137 -88 -13131 88
rect -13097 -88 -13091 88
rect -13137 -100 -13091 -88
rect -12979 88 -12933 100
rect -12979 -88 -12973 88
rect -12939 -88 -12933 88
rect -12979 -100 -12933 -88
rect -12821 88 -12775 100
rect -12821 -88 -12815 88
rect -12781 -88 -12775 88
rect -12821 -100 -12775 -88
rect -12663 88 -12617 100
rect -12663 -88 -12657 88
rect -12623 -88 -12617 88
rect -12663 -100 -12617 -88
rect -12505 88 -12459 100
rect -12505 -88 -12499 88
rect -12465 -88 -12459 88
rect -12505 -100 -12459 -88
rect -12347 88 -12301 100
rect -12347 -88 -12341 88
rect -12307 -88 -12301 88
rect -12347 -100 -12301 -88
rect -12189 88 -12143 100
rect -12189 -88 -12183 88
rect -12149 -88 -12143 88
rect -12189 -100 -12143 -88
rect -12031 88 -11985 100
rect -12031 -88 -12025 88
rect -11991 -88 -11985 88
rect -12031 -100 -11985 -88
rect -11873 88 -11827 100
rect -11873 -88 -11867 88
rect -11833 -88 -11827 88
rect -11873 -100 -11827 -88
rect -11715 88 -11669 100
rect -11715 -88 -11709 88
rect -11675 -88 -11669 88
rect -11715 -100 -11669 -88
rect -11557 88 -11511 100
rect -11557 -88 -11551 88
rect -11517 -88 -11511 88
rect -11557 -100 -11511 -88
rect -11399 88 -11353 100
rect -11399 -88 -11393 88
rect -11359 -88 -11353 88
rect -11399 -100 -11353 -88
rect -11241 88 -11195 100
rect -11241 -88 -11235 88
rect -11201 -88 -11195 88
rect -11241 -100 -11195 -88
rect -11083 88 -11037 100
rect -11083 -88 -11077 88
rect -11043 -88 -11037 88
rect -11083 -100 -11037 -88
rect -10925 88 -10879 100
rect -10925 -88 -10919 88
rect -10885 -88 -10879 88
rect -10925 -100 -10879 -88
rect -10767 88 -10721 100
rect -10767 -88 -10761 88
rect -10727 -88 -10721 88
rect -10767 -100 -10721 -88
rect -10609 88 -10563 100
rect -10609 -88 -10603 88
rect -10569 -88 -10563 88
rect -10609 -100 -10563 -88
rect -10451 88 -10405 100
rect -10451 -88 -10445 88
rect -10411 -88 -10405 88
rect -10451 -100 -10405 -88
rect -10293 88 -10247 100
rect -10293 -88 -10287 88
rect -10253 -88 -10247 88
rect -10293 -100 -10247 -88
rect -10135 88 -10089 100
rect -10135 -88 -10129 88
rect -10095 -88 -10089 88
rect -10135 -100 -10089 -88
rect -9977 88 -9931 100
rect -9977 -88 -9971 88
rect -9937 -88 -9931 88
rect -9977 -100 -9931 -88
rect -9819 88 -9773 100
rect -9819 -88 -9813 88
rect -9779 -88 -9773 88
rect -9819 -100 -9773 -88
rect -9661 88 -9615 100
rect -9661 -88 -9655 88
rect -9621 -88 -9615 88
rect -9661 -100 -9615 -88
rect -9503 88 -9457 100
rect -9503 -88 -9497 88
rect -9463 -88 -9457 88
rect -9503 -100 -9457 -88
rect -9345 88 -9299 100
rect -9345 -88 -9339 88
rect -9305 -88 -9299 88
rect -9345 -100 -9299 -88
rect -9187 88 -9141 100
rect -9187 -88 -9181 88
rect -9147 -88 -9141 88
rect -9187 -100 -9141 -88
rect -9029 88 -8983 100
rect -9029 -88 -9023 88
rect -8989 -88 -8983 88
rect -9029 -100 -8983 -88
rect -8871 88 -8825 100
rect -8871 -88 -8865 88
rect -8831 -88 -8825 88
rect -8871 -100 -8825 -88
rect -8713 88 -8667 100
rect -8713 -88 -8707 88
rect -8673 -88 -8667 88
rect -8713 -100 -8667 -88
rect -8555 88 -8509 100
rect -8555 -88 -8549 88
rect -8515 -88 -8509 88
rect -8555 -100 -8509 -88
rect -8397 88 -8351 100
rect -8397 -88 -8391 88
rect -8357 -88 -8351 88
rect -8397 -100 -8351 -88
rect -8239 88 -8193 100
rect -8239 -88 -8233 88
rect -8199 -88 -8193 88
rect -8239 -100 -8193 -88
rect -8081 88 -8035 100
rect -8081 -88 -8075 88
rect -8041 -88 -8035 88
rect -8081 -100 -8035 -88
rect -7923 88 -7877 100
rect -7923 -88 -7917 88
rect -7883 -88 -7877 88
rect -7923 -100 -7877 -88
rect -7765 88 -7719 100
rect -7765 -88 -7759 88
rect -7725 -88 -7719 88
rect -7765 -100 -7719 -88
rect -7607 88 -7561 100
rect -7607 -88 -7601 88
rect -7567 -88 -7561 88
rect -7607 -100 -7561 -88
rect -7449 88 -7403 100
rect -7449 -88 -7443 88
rect -7409 -88 -7403 88
rect -7449 -100 -7403 -88
rect -7291 88 -7245 100
rect -7291 -88 -7285 88
rect -7251 -88 -7245 88
rect -7291 -100 -7245 -88
rect -7133 88 -7087 100
rect -7133 -88 -7127 88
rect -7093 -88 -7087 88
rect -7133 -100 -7087 -88
rect -6975 88 -6929 100
rect -6975 -88 -6969 88
rect -6935 -88 -6929 88
rect -6975 -100 -6929 -88
rect -6817 88 -6771 100
rect -6817 -88 -6811 88
rect -6777 -88 -6771 88
rect -6817 -100 -6771 -88
rect -6659 88 -6613 100
rect -6659 -88 -6653 88
rect -6619 -88 -6613 88
rect -6659 -100 -6613 -88
rect -6501 88 -6455 100
rect -6501 -88 -6495 88
rect -6461 -88 -6455 88
rect -6501 -100 -6455 -88
rect -6343 88 -6297 100
rect -6343 -88 -6337 88
rect -6303 -88 -6297 88
rect -6343 -100 -6297 -88
rect -6185 88 -6139 100
rect -6185 -88 -6179 88
rect -6145 -88 -6139 88
rect -6185 -100 -6139 -88
rect -6027 88 -5981 100
rect -6027 -88 -6021 88
rect -5987 -88 -5981 88
rect -6027 -100 -5981 -88
rect -5869 88 -5823 100
rect -5869 -88 -5863 88
rect -5829 -88 -5823 88
rect -5869 -100 -5823 -88
rect -5711 88 -5665 100
rect -5711 -88 -5705 88
rect -5671 -88 -5665 88
rect -5711 -100 -5665 -88
rect -5553 88 -5507 100
rect -5553 -88 -5547 88
rect -5513 -88 -5507 88
rect -5553 -100 -5507 -88
rect -5395 88 -5349 100
rect -5395 -88 -5389 88
rect -5355 -88 -5349 88
rect -5395 -100 -5349 -88
rect -5237 88 -5191 100
rect -5237 -88 -5231 88
rect -5197 -88 -5191 88
rect -5237 -100 -5191 -88
rect -5079 88 -5033 100
rect -5079 -88 -5073 88
rect -5039 -88 -5033 88
rect -5079 -100 -5033 -88
rect -4921 88 -4875 100
rect -4921 -88 -4915 88
rect -4881 -88 -4875 88
rect -4921 -100 -4875 -88
rect -4763 88 -4717 100
rect -4763 -88 -4757 88
rect -4723 -88 -4717 88
rect -4763 -100 -4717 -88
rect -4605 88 -4559 100
rect -4605 -88 -4599 88
rect -4565 -88 -4559 88
rect -4605 -100 -4559 -88
rect -4447 88 -4401 100
rect -4447 -88 -4441 88
rect -4407 -88 -4401 88
rect -4447 -100 -4401 -88
rect -4289 88 -4243 100
rect -4289 -88 -4283 88
rect -4249 -88 -4243 88
rect -4289 -100 -4243 -88
rect -4131 88 -4085 100
rect -4131 -88 -4125 88
rect -4091 -88 -4085 88
rect -4131 -100 -4085 -88
rect -3973 88 -3927 100
rect -3973 -88 -3967 88
rect -3933 -88 -3927 88
rect -3973 -100 -3927 -88
rect -3815 88 -3769 100
rect -3815 -88 -3809 88
rect -3775 -88 -3769 88
rect -3815 -100 -3769 -88
rect -3657 88 -3611 100
rect -3657 -88 -3651 88
rect -3617 -88 -3611 88
rect -3657 -100 -3611 -88
rect -3499 88 -3453 100
rect -3499 -88 -3493 88
rect -3459 -88 -3453 88
rect -3499 -100 -3453 -88
rect -3341 88 -3295 100
rect -3341 -88 -3335 88
rect -3301 -88 -3295 88
rect -3341 -100 -3295 -88
rect -3183 88 -3137 100
rect -3183 -88 -3177 88
rect -3143 -88 -3137 88
rect -3183 -100 -3137 -88
rect -3025 88 -2979 100
rect -3025 -88 -3019 88
rect -2985 -88 -2979 88
rect -3025 -100 -2979 -88
rect -2867 88 -2821 100
rect -2867 -88 -2861 88
rect -2827 -88 -2821 88
rect -2867 -100 -2821 -88
rect -2709 88 -2663 100
rect -2709 -88 -2703 88
rect -2669 -88 -2663 88
rect -2709 -100 -2663 -88
rect -2551 88 -2505 100
rect -2551 -88 -2545 88
rect -2511 -88 -2505 88
rect -2551 -100 -2505 -88
rect -2393 88 -2347 100
rect -2393 -88 -2387 88
rect -2353 -88 -2347 88
rect -2393 -100 -2347 -88
rect -2235 88 -2189 100
rect -2235 -88 -2229 88
rect -2195 -88 -2189 88
rect -2235 -100 -2189 -88
rect -2077 88 -2031 100
rect -2077 -88 -2071 88
rect -2037 -88 -2031 88
rect -2077 -100 -2031 -88
rect -1919 88 -1873 100
rect -1919 -88 -1913 88
rect -1879 -88 -1873 88
rect -1919 -100 -1873 -88
rect -1761 88 -1715 100
rect -1761 -88 -1755 88
rect -1721 -88 -1715 88
rect -1761 -100 -1715 -88
rect -1603 88 -1557 100
rect -1603 -88 -1597 88
rect -1563 -88 -1557 88
rect -1603 -100 -1557 -88
rect -1445 88 -1399 100
rect -1445 -88 -1439 88
rect -1405 -88 -1399 88
rect -1445 -100 -1399 -88
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect 1399 88 1445 100
rect 1399 -88 1405 88
rect 1439 -88 1445 88
rect 1399 -100 1445 -88
rect 1557 88 1603 100
rect 1557 -88 1563 88
rect 1597 -88 1603 88
rect 1557 -100 1603 -88
rect 1715 88 1761 100
rect 1715 -88 1721 88
rect 1755 -88 1761 88
rect 1715 -100 1761 -88
rect 1873 88 1919 100
rect 1873 -88 1879 88
rect 1913 -88 1919 88
rect 1873 -100 1919 -88
rect 2031 88 2077 100
rect 2031 -88 2037 88
rect 2071 -88 2077 88
rect 2031 -100 2077 -88
rect 2189 88 2235 100
rect 2189 -88 2195 88
rect 2229 -88 2235 88
rect 2189 -100 2235 -88
rect 2347 88 2393 100
rect 2347 -88 2353 88
rect 2387 -88 2393 88
rect 2347 -100 2393 -88
rect 2505 88 2551 100
rect 2505 -88 2511 88
rect 2545 -88 2551 88
rect 2505 -100 2551 -88
rect 2663 88 2709 100
rect 2663 -88 2669 88
rect 2703 -88 2709 88
rect 2663 -100 2709 -88
rect 2821 88 2867 100
rect 2821 -88 2827 88
rect 2861 -88 2867 88
rect 2821 -100 2867 -88
rect 2979 88 3025 100
rect 2979 -88 2985 88
rect 3019 -88 3025 88
rect 2979 -100 3025 -88
rect 3137 88 3183 100
rect 3137 -88 3143 88
rect 3177 -88 3183 88
rect 3137 -100 3183 -88
rect 3295 88 3341 100
rect 3295 -88 3301 88
rect 3335 -88 3341 88
rect 3295 -100 3341 -88
rect 3453 88 3499 100
rect 3453 -88 3459 88
rect 3493 -88 3499 88
rect 3453 -100 3499 -88
rect 3611 88 3657 100
rect 3611 -88 3617 88
rect 3651 -88 3657 88
rect 3611 -100 3657 -88
rect 3769 88 3815 100
rect 3769 -88 3775 88
rect 3809 -88 3815 88
rect 3769 -100 3815 -88
rect 3927 88 3973 100
rect 3927 -88 3933 88
rect 3967 -88 3973 88
rect 3927 -100 3973 -88
rect 4085 88 4131 100
rect 4085 -88 4091 88
rect 4125 -88 4131 88
rect 4085 -100 4131 -88
rect 4243 88 4289 100
rect 4243 -88 4249 88
rect 4283 -88 4289 88
rect 4243 -100 4289 -88
rect 4401 88 4447 100
rect 4401 -88 4407 88
rect 4441 -88 4447 88
rect 4401 -100 4447 -88
rect 4559 88 4605 100
rect 4559 -88 4565 88
rect 4599 -88 4605 88
rect 4559 -100 4605 -88
rect 4717 88 4763 100
rect 4717 -88 4723 88
rect 4757 -88 4763 88
rect 4717 -100 4763 -88
rect 4875 88 4921 100
rect 4875 -88 4881 88
rect 4915 -88 4921 88
rect 4875 -100 4921 -88
rect 5033 88 5079 100
rect 5033 -88 5039 88
rect 5073 -88 5079 88
rect 5033 -100 5079 -88
rect 5191 88 5237 100
rect 5191 -88 5197 88
rect 5231 -88 5237 88
rect 5191 -100 5237 -88
rect 5349 88 5395 100
rect 5349 -88 5355 88
rect 5389 -88 5395 88
rect 5349 -100 5395 -88
rect 5507 88 5553 100
rect 5507 -88 5513 88
rect 5547 -88 5553 88
rect 5507 -100 5553 -88
rect 5665 88 5711 100
rect 5665 -88 5671 88
rect 5705 -88 5711 88
rect 5665 -100 5711 -88
rect 5823 88 5869 100
rect 5823 -88 5829 88
rect 5863 -88 5869 88
rect 5823 -100 5869 -88
rect 5981 88 6027 100
rect 5981 -88 5987 88
rect 6021 -88 6027 88
rect 5981 -100 6027 -88
rect 6139 88 6185 100
rect 6139 -88 6145 88
rect 6179 -88 6185 88
rect 6139 -100 6185 -88
rect 6297 88 6343 100
rect 6297 -88 6303 88
rect 6337 -88 6343 88
rect 6297 -100 6343 -88
rect 6455 88 6501 100
rect 6455 -88 6461 88
rect 6495 -88 6501 88
rect 6455 -100 6501 -88
rect 6613 88 6659 100
rect 6613 -88 6619 88
rect 6653 -88 6659 88
rect 6613 -100 6659 -88
rect 6771 88 6817 100
rect 6771 -88 6777 88
rect 6811 -88 6817 88
rect 6771 -100 6817 -88
rect 6929 88 6975 100
rect 6929 -88 6935 88
rect 6969 -88 6975 88
rect 6929 -100 6975 -88
rect 7087 88 7133 100
rect 7087 -88 7093 88
rect 7127 -88 7133 88
rect 7087 -100 7133 -88
rect 7245 88 7291 100
rect 7245 -88 7251 88
rect 7285 -88 7291 88
rect 7245 -100 7291 -88
rect 7403 88 7449 100
rect 7403 -88 7409 88
rect 7443 -88 7449 88
rect 7403 -100 7449 -88
rect 7561 88 7607 100
rect 7561 -88 7567 88
rect 7601 -88 7607 88
rect 7561 -100 7607 -88
rect 7719 88 7765 100
rect 7719 -88 7725 88
rect 7759 -88 7765 88
rect 7719 -100 7765 -88
rect 7877 88 7923 100
rect 7877 -88 7883 88
rect 7917 -88 7923 88
rect 7877 -100 7923 -88
rect 8035 88 8081 100
rect 8035 -88 8041 88
rect 8075 -88 8081 88
rect 8035 -100 8081 -88
rect 8193 88 8239 100
rect 8193 -88 8199 88
rect 8233 -88 8239 88
rect 8193 -100 8239 -88
rect 8351 88 8397 100
rect 8351 -88 8357 88
rect 8391 -88 8397 88
rect 8351 -100 8397 -88
rect 8509 88 8555 100
rect 8509 -88 8515 88
rect 8549 -88 8555 88
rect 8509 -100 8555 -88
rect 8667 88 8713 100
rect 8667 -88 8673 88
rect 8707 -88 8713 88
rect 8667 -100 8713 -88
rect 8825 88 8871 100
rect 8825 -88 8831 88
rect 8865 -88 8871 88
rect 8825 -100 8871 -88
rect 8983 88 9029 100
rect 8983 -88 8989 88
rect 9023 -88 9029 88
rect 8983 -100 9029 -88
rect 9141 88 9187 100
rect 9141 -88 9147 88
rect 9181 -88 9187 88
rect 9141 -100 9187 -88
rect 9299 88 9345 100
rect 9299 -88 9305 88
rect 9339 -88 9345 88
rect 9299 -100 9345 -88
rect 9457 88 9503 100
rect 9457 -88 9463 88
rect 9497 -88 9503 88
rect 9457 -100 9503 -88
rect 9615 88 9661 100
rect 9615 -88 9621 88
rect 9655 -88 9661 88
rect 9615 -100 9661 -88
rect 9773 88 9819 100
rect 9773 -88 9779 88
rect 9813 -88 9819 88
rect 9773 -100 9819 -88
rect 9931 88 9977 100
rect 9931 -88 9937 88
rect 9971 -88 9977 88
rect 9931 -100 9977 -88
rect 10089 88 10135 100
rect 10089 -88 10095 88
rect 10129 -88 10135 88
rect 10089 -100 10135 -88
rect 10247 88 10293 100
rect 10247 -88 10253 88
rect 10287 -88 10293 88
rect 10247 -100 10293 -88
rect 10405 88 10451 100
rect 10405 -88 10411 88
rect 10445 -88 10451 88
rect 10405 -100 10451 -88
rect 10563 88 10609 100
rect 10563 -88 10569 88
rect 10603 -88 10609 88
rect 10563 -100 10609 -88
rect 10721 88 10767 100
rect 10721 -88 10727 88
rect 10761 -88 10767 88
rect 10721 -100 10767 -88
rect 10879 88 10925 100
rect 10879 -88 10885 88
rect 10919 -88 10925 88
rect 10879 -100 10925 -88
rect 11037 88 11083 100
rect 11037 -88 11043 88
rect 11077 -88 11083 88
rect 11037 -100 11083 -88
rect 11195 88 11241 100
rect 11195 -88 11201 88
rect 11235 -88 11241 88
rect 11195 -100 11241 -88
rect 11353 88 11399 100
rect 11353 -88 11359 88
rect 11393 -88 11399 88
rect 11353 -100 11399 -88
rect 11511 88 11557 100
rect 11511 -88 11517 88
rect 11551 -88 11557 88
rect 11511 -100 11557 -88
rect 11669 88 11715 100
rect 11669 -88 11675 88
rect 11709 -88 11715 88
rect 11669 -100 11715 -88
rect 11827 88 11873 100
rect 11827 -88 11833 88
rect 11867 -88 11873 88
rect 11827 -100 11873 -88
rect 11985 88 12031 100
rect 11985 -88 11991 88
rect 12025 -88 12031 88
rect 11985 -100 12031 -88
rect 12143 88 12189 100
rect 12143 -88 12149 88
rect 12183 -88 12189 88
rect 12143 -100 12189 -88
rect 12301 88 12347 100
rect 12301 -88 12307 88
rect 12341 -88 12347 88
rect 12301 -100 12347 -88
rect 12459 88 12505 100
rect 12459 -88 12465 88
rect 12499 -88 12505 88
rect 12459 -100 12505 -88
rect 12617 88 12663 100
rect 12617 -88 12623 88
rect 12657 -88 12663 88
rect 12617 -100 12663 -88
rect 12775 88 12821 100
rect 12775 -88 12781 88
rect 12815 -88 12821 88
rect 12775 -100 12821 -88
rect 12933 88 12979 100
rect 12933 -88 12939 88
rect 12973 -88 12979 88
rect 12933 -100 12979 -88
rect 13091 88 13137 100
rect 13091 -88 13097 88
rect 13131 -88 13137 88
rect 13091 -100 13137 -88
rect 13249 88 13295 100
rect 13249 -88 13255 88
rect 13289 -88 13295 88
rect 13249 -100 13295 -88
rect 13407 88 13453 100
rect 13407 -88 13413 88
rect 13447 -88 13453 88
rect 13407 -100 13453 -88
rect 13565 88 13611 100
rect 13565 -88 13571 88
rect 13605 -88 13611 88
rect 13565 -100 13611 -88
rect 13723 88 13769 100
rect 13723 -88 13729 88
rect 13763 -88 13769 88
rect 13723 -100 13769 -88
rect 13881 88 13927 100
rect 13881 -88 13887 88
rect 13921 -88 13927 88
rect 13881 -100 13927 -88
rect 14039 88 14085 100
rect 14039 -88 14045 88
rect 14079 -88 14085 88
rect 14039 -100 14085 -88
rect 14197 88 14243 100
rect 14197 -88 14203 88
rect 14237 -88 14243 88
rect 14197 -100 14243 -88
rect 14355 88 14401 100
rect 14355 -88 14361 88
rect 14395 -88 14401 88
rect 14355 -100 14401 -88
rect 14513 88 14559 100
rect 14513 -88 14519 88
rect 14553 -88 14559 88
rect 14513 -100 14559 -88
rect 14671 88 14717 100
rect 14671 -88 14677 88
rect 14711 -88 14717 88
rect 14671 -100 14717 -88
rect 14829 88 14875 100
rect 14829 -88 14835 88
rect 14869 -88 14875 88
rect 14829 -100 14875 -88
rect 14987 88 15033 100
rect 14987 -88 14993 88
rect 15027 -88 15033 88
rect 14987 -100 15033 -88
rect 15145 88 15191 100
rect 15145 -88 15151 88
rect 15185 -88 15191 88
rect 15145 -100 15191 -88
rect 15303 88 15349 100
rect 15303 -88 15309 88
rect 15343 -88 15349 88
rect 15303 -100 15349 -88
rect 15461 88 15507 100
rect 15461 -88 15467 88
rect 15501 -88 15507 88
rect 15461 -100 15507 -88
rect 15619 88 15665 100
rect 15619 -88 15625 88
rect 15659 -88 15665 88
rect 15619 -100 15665 -88
rect 15777 88 15823 100
rect 15777 -88 15783 88
rect 15817 -88 15823 88
rect 15777 -100 15823 -88
rect -15767 -147 -15675 -141
rect -15767 -181 -15755 -147
rect -15687 -181 -15675 -147
rect -15767 -187 -15675 -181
rect -15609 -147 -15517 -141
rect -15609 -181 -15597 -147
rect -15529 -181 -15517 -147
rect -15609 -187 -15517 -181
rect -15451 -147 -15359 -141
rect -15451 -181 -15439 -147
rect -15371 -181 -15359 -147
rect -15451 -187 -15359 -181
rect -15293 -147 -15201 -141
rect -15293 -181 -15281 -147
rect -15213 -181 -15201 -147
rect -15293 -187 -15201 -181
rect -15135 -147 -15043 -141
rect -15135 -181 -15123 -147
rect -15055 -181 -15043 -147
rect -15135 -187 -15043 -181
rect -14977 -147 -14885 -141
rect -14977 -181 -14965 -147
rect -14897 -181 -14885 -147
rect -14977 -187 -14885 -181
rect -14819 -147 -14727 -141
rect -14819 -181 -14807 -147
rect -14739 -181 -14727 -147
rect -14819 -187 -14727 -181
rect -14661 -147 -14569 -141
rect -14661 -181 -14649 -147
rect -14581 -181 -14569 -147
rect -14661 -187 -14569 -181
rect -14503 -147 -14411 -141
rect -14503 -181 -14491 -147
rect -14423 -181 -14411 -147
rect -14503 -187 -14411 -181
rect -14345 -147 -14253 -141
rect -14345 -181 -14333 -147
rect -14265 -181 -14253 -147
rect -14345 -187 -14253 -181
rect -14187 -147 -14095 -141
rect -14187 -181 -14175 -147
rect -14107 -181 -14095 -147
rect -14187 -187 -14095 -181
rect -14029 -147 -13937 -141
rect -14029 -181 -14017 -147
rect -13949 -181 -13937 -147
rect -14029 -187 -13937 -181
rect -13871 -147 -13779 -141
rect -13871 -181 -13859 -147
rect -13791 -181 -13779 -147
rect -13871 -187 -13779 -181
rect -13713 -147 -13621 -141
rect -13713 -181 -13701 -147
rect -13633 -181 -13621 -147
rect -13713 -187 -13621 -181
rect -13555 -147 -13463 -141
rect -13555 -181 -13543 -147
rect -13475 -181 -13463 -147
rect -13555 -187 -13463 -181
rect -13397 -147 -13305 -141
rect -13397 -181 -13385 -147
rect -13317 -181 -13305 -147
rect -13397 -187 -13305 -181
rect -13239 -147 -13147 -141
rect -13239 -181 -13227 -147
rect -13159 -181 -13147 -147
rect -13239 -187 -13147 -181
rect -13081 -147 -12989 -141
rect -13081 -181 -13069 -147
rect -13001 -181 -12989 -147
rect -13081 -187 -12989 -181
rect -12923 -147 -12831 -141
rect -12923 -181 -12911 -147
rect -12843 -181 -12831 -147
rect -12923 -187 -12831 -181
rect -12765 -147 -12673 -141
rect -12765 -181 -12753 -147
rect -12685 -181 -12673 -147
rect -12765 -187 -12673 -181
rect -12607 -147 -12515 -141
rect -12607 -181 -12595 -147
rect -12527 -181 -12515 -147
rect -12607 -187 -12515 -181
rect -12449 -147 -12357 -141
rect -12449 -181 -12437 -147
rect -12369 -181 -12357 -147
rect -12449 -187 -12357 -181
rect -12291 -147 -12199 -141
rect -12291 -181 -12279 -147
rect -12211 -181 -12199 -147
rect -12291 -187 -12199 -181
rect -12133 -147 -12041 -141
rect -12133 -181 -12121 -147
rect -12053 -181 -12041 -147
rect -12133 -187 -12041 -181
rect -11975 -147 -11883 -141
rect -11975 -181 -11963 -147
rect -11895 -181 -11883 -147
rect -11975 -187 -11883 -181
rect -11817 -147 -11725 -141
rect -11817 -181 -11805 -147
rect -11737 -181 -11725 -147
rect -11817 -187 -11725 -181
rect -11659 -147 -11567 -141
rect -11659 -181 -11647 -147
rect -11579 -181 -11567 -147
rect -11659 -187 -11567 -181
rect -11501 -147 -11409 -141
rect -11501 -181 -11489 -147
rect -11421 -181 -11409 -147
rect -11501 -187 -11409 -181
rect -11343 -147 -11251 -141
rect -11343 -181 -11331 -147
rect -11263 -181 -11251 -147
rect -11343 -187 -11251 -181
rect -11185 -147 -11093 -141
rect -11185 -181 -11173 -147
rect -11105 -181 -11093 -147
rect -11185 -187 -11093 -181
rect -11027 -147 -10935 -141
rect -11027 -181 -11015 -147
rect -10947 -181 -10935 -147
rect -11027 -187 -10935 -181
rect -10869 -147 -10777 -141
rect -10869 -181 -10857 -147
rect -10789 -181 -10777 -147
rect -10869 -187 -10777 -181
rect -10711 -147 -10619 -141
rect -10711 -181 -10699 -147
rect -10631 -181 -10619 -147
rect -10711 -187 -10619 -181
rect -10553 -147 -10461 -141
rect -10553 -181 -10541 -147
rect -10473 -181 -10461 -147
rect -10553 -187 -10461 -181
rect -10395 -147 -10303 -141
rect -10395 -181 -10383 -147
rect -10315 -181 -10303 -147
rect -10395 -187 -10303 -181
rect -10237 -147 -10145 -141
rect -10237 -181 -10225 -147
rect -10157 -181 -10145 -147
rect -10237 -187 -10145 -181
rect -10079 -147 -9987 -141
rect -10079 -181 -10067 -147
rect -9999 -181 -9987 -147
rect -10079 -187 -9987 -181
rect -9921 -147 -9829 -141
rect -9921 -181 -9909 -147
rect -9841 -181 -9829 -147
rect -9921 -187 -9829 -181
rect -9763 -147 -9671 -141
rect -9763 -181 -9751 -147
rect -9683 -181 -9671 -147
rect -9763 -187 -9671 -181
rect -9605 -147 -9513 -141
rect -9605 -181 -9593 -147
rect -9525 -181 -9513 -147
rect -9605 -187 -9513 -181
rect -9447 -147 -9355 -141
rect -9447 -181 -9435 -147
rect -9367 -181 -9355 -147
rect -9447 -187 -9355 -181
rect -9289 -147 -9197 -141
rect -9289 -181 -9277 -147
rect -9209 -181 -9197 -147
rect -9289 -187 -9197 -181
rect -9131 -147 -9039 -141
rect -9131 -181 -9119 -147
rect -9051 -181 -9039 -147
rect -9131 -187 -9039 -181
rect -8973 -147 -8881 -141
rect -8973 -181 -8961 -147
rect -8893 -181 -8881 -147
rect -8973 -187 -8881 -181
rect -8815 -147 -8723 -141
rect -8815 -181 -8803 -147
rect -8735 -181 -8723 -147
rect -8815 -187 -8723 -181
rect -8657 -147 -8565 -141
rect -8657 -181 -8645 -147
rect -8577 -181 -8565 -147
rect -8657 -187 -8565 -181
rect -8499 -147 -8407 -141
rect -8499 -181 -8487 -147
rect -8419 -181 -8407 -147
rect -8499 -187 -8407 -181
rect -8341 -147 -8249 -141
rect -8341 -181 -8329 -147
rect -8261 -181 -8249 -147
rect -8341 -187 -8249 -181
rect -8183 -147 -8091 -141
rect -8183 -181 -8171 -147
rect -8103 -181 -8091 -147
rect -8183 -187 -8091 -181
rect -8025 -147 -7933 -141
rect -8025 -181 -8013 -147
rect -7945 -181 -7933 -147
rect -8025 -187 -7933 -181
rect -7867 -147 -7775 -141
rect -7867 -181 -7855 -147
rect -7787 -181 -7775 -147
rect -7867 -187 -7775 -181
rect -7709 -147 -7617 -141
rect -7709 -181 -7697 -147
rect -7629 -181 -7617 -147
rect -7709 -187 -7617 -181
rect -7551 -147 -7459 -141
rect -7551 -181 -7539 -147
rect -7471 -181 -7459 -147
rect -7551 -187 -7459 -181
rect -7393 -147 -7301 -141
rect -7393 -181 -7381 -147
rect -7313 -181 -7301 -147
rect -7393 -187 -7301 -181
rect -7235 -147 -7143 -141
rect -7235 -181 -7223 -147
rect -7155 -181 -7143 -147
rect -7235 -187 -7143 -181
rect -7077 -147 -6985 -141
rect -7077 -181 -7065 -147
rect -6997 -181 -6985 -147
rect -7077 -187 -6985 -181
rect -6919 -147 -6827 -141
rect -6919 -181 -6907 -147
rect -6839 -181 -6827 -147
rect -6919 -187 -6827 -181
rect -6761 -147 -6669 -141
rect -6761 -181 -6749 -147
rect -6681 -181 -6669 -147
rect -6761 -187 -6669 -181
rect -6603 -147 -6511 -141
rect -6603 -181 -6591 -147
rect -6523 -181 -6511 -147
rect -6603 -187 -6511 -181
rect -6445 -147 -6353 -141
rect -6445 -181 -6433 -147
rect -6365 -181 -6353 -147
rect -6445 -187 -6353 -181
rect -6287 -147 -6195 -141
rect -6287 -181 -6275 -147
rect -6207 -181 -6195 -147
rect -6287 -187 -6195 -181
rect -6129 -147 -6037 -141
rect -6129 -181 -6117 -147
rect -6049 -181 -6037 -147
rect -6129 -187 -6037 -181
rect -5971 -147 -5879 -141
rect -5971 -181 -5959 -147
rect -5891 -181 -5879 -147
rect -5971 -187 -5879 -181
rect -5813 -147 -5721 -141
rect -5813 -181 -5801 -147
rect -5733 -181 -5721 -147
rect -5813 -187 -5721 -181
rect -5655 -147 -5563 -141
rect -5655 -181 -5643 -147
rect -5575 -181 -5563 -147
rect -5655 -187 -5563 -181
rect -5497 -147 -5405 -141
rect -5497 -181 -5485 -147
rect -5417 -181 -5405 -147
rect -5497 -187 -5405 -181
rect -5339 -147 -5247 -141
rect -5339 -181 -5327 -147
rect -5259 -181 -5247 -147
rect -5339 -187 -5247 -181
rect -5181 -147 -5089 -141
rect -5181 -181 -5169 -147
rect -5101 -181 -5089 -147
rect -5181 -187 -5089 -181
rect -5023 -147 -4931 -141
rect -5023 -181 -5011 -147
rect -4943 -181 -4931 -147
rect -5023 -187 -4931 -181
rect -4865 -147 -4773 -141
rect -4865 -181 -4853 -147
rect -4785 -181 -4773 -147
rect -4865 -187 -4773 -181
rect -4707 -147 -4615 -141
rect -4707 -181 -4695 -147
rect -4627 -181 -4615 -147
rect -4707 -187 -4615 -181
rect -4549 -147 -4457 -141
rect -4549 -181 -4537 -147
rect -4469 -181 -4457 -147
rect -4549 -187 -4457 -181
rect -4391 -147 -4299 -141
rect -4391 -181 -4379 -147
rect -4311 -181 -4299 -147
rect -4391 -187 -4299 -181
rect -4233 -147 -4141 -141
rect -4233 -181 -4221 -147
rect -4153 -181 -4141 -147
rect -4233 -187 -4141 -181
rect -4075 -147 -3983 -141
rect -4075 -181 -4063 -147
rect -3995 -181 -3983 -147
rect -4075 -187 -3983 -181
rect -3917 -147 -3825 -141
rect -3917 -181 -3905 -147
rect -3837 -181 -3825 -147
rect -3917 -187 -3825 -181
rect -3759 -147 -3667 -141
rect -3759 -181 -3747 -147
rect -3679 -181 -3667 -147
rect -3759 -187 -3667 -181
rect -3601 -147 -3509 -141
rect -3601 -181 -3589 -147
rect -3521 -181 -3509 -147
rect -3601 -187 -3509 -181
rect -3443 -147 -3351 -141
rect -3443 -181 -3431 -147
rect -3363 -181 -3351 -147
rect -3443 -187 -3351 -181
rect -3285 -147 -3193 -141
rect -3285 -181 -3273 -147
rect -3205 -181 -3193 -147
rect -3285 -187 -3193 -181
rect -3127 -147 -3035 -141
rect -3127 -181 -3115 -147
rect -3047 -181 -3035 -147
rect -3127 -187 -3035 -181
rect -2969 -147 -2877 -141
rect -2969 -181 -2957 -147
rect -2889 -181 -2877 -147
rect -2969 -187 -2877 -181
rect -2811 -147 -2719 -141
rect -2811 -181 -2799 -147
rect -2731 -181 -2719 -147
rect -2811 -187 -2719 -181
rect -2653 -147 -2561 -141
rect -2653 -181 -2641 -147
rect -2573 -181 -2561 -147
rect -2653 -187 -2561 -181
rect -2495 -147 -2403 -141
rect -2495 -181 -2483 -147
rect -2415 -181 -2403 -147
rect -2495 -187 -2403 -181
rect -2337 -147 -2245 -141
rect -2337 -181 -2325 -147
rect -2257 -181 -2245 -147
rect -2337 -187 -2245 -181
rect -2179 -147 -2087 -141
rect -2179 -181 -2167 -147
rect -2099 -181 -2087 -147
rect -2179 -187 -2087 -181
rect -2021 -147 -1929 -141
rect -2021 -181 -2009 -147
rect -1941 -181 -1929 -147
rect -2021 -187 -1929 -181
rect -1863 -147 -1771 -141
rect -1863 -181 -1851 -147
rect -1783 -181 -1771 -147
rect -1863 -187 -1771 -181
rect -1705 -147 -1613 -141
rect -1705 -181 -1693 -147
rect -1625 -181 -1613 -147
rect -1705 -187 -1613 -181
rect -1547 -147 -1455 -141
rect -1547 -181 -1535 -147
rect -1467 -181 -1455 -147
rect -1547 -187 -1455 -181
rect -1389 -147 -1297 -141
rect -1389 -181 -1377 -147
rect -1309 -181 -1297 -147
rect -1389 -187 -1297 -181
rect -1231 -147 -1139 -141
rect -1231 -181 -1219 -147
rect -1151 -181 -1139 -147
rect -1231 -187 -1139 -181
rect -1073 -147 -981 -141
rect -1073 -181 -1061 -147
rect -993 -181 -981 -147
rect -1073 -187 -981 -181
rect -915 -147 -823 -141
rect -915 -181 -903 -147
rect -835 -181 -823 -147
rect -915 -187 -823 -181
rect -757 -147 -665 -141
rect -757 -181 -745 -147
rect -677 -181 -665 -147
rect -757 -187 -665 -181
rect -599 -147 -507 -141
rect -599 -181 -587 -147
rect -519 -181 -507 -147
rect -599 -187 -507 -181
rect -441 -147 -349 -141
rect -441 -181 -429 -147
rect -361 -181 -349 -147
rect -441 -187 -349 -181
rect -283 -147 -191 -141
rect -283 -181 -271 -147
rect -203 -181 -191 -147
rect -283 -187 -191 -181
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
rect 191 -147 283 -141
rect 191 -181 203 -147
rect 271 -181 283 -147
rect 191 -187 283 -181
rect 349 -147 441 -141
rect 349 -181 361 -147
rect 429 -181 441 -147
rect 349 -187 441 -181
rect 507 -147 599 -141
rect 507 -181 519 -147
rect 587 -181 599 -147
rect 507 -187 599 -181
rect 665 -147 757 -141
rect 665 -181 677 -147
rect 745 -181 757 -147
rect 665 -187 757 -181
rect 823 -147 915 -141
rect 823 -181 835 -147
rect 903 -181 915 -147
rect 823 -187 915 -181
rect 981 -147 1073 -141
rect 981 -181 993 -147
rect 1061 -181 1073 -147
rect 981 -187 1073 -181
rect 1139 -147 1231 -141
rect 1139 -181 1151 -147
rect 1219 -181 1231 -147
rect 1139 -187 1231 -181
rect 1297 -147 1389 -141
rect 1297 -181 1309 -147
rect 1377 -181 1389 -147
rect 1297 -187 1389 -181
rect 1455 -147 1547 -141
rect 1455 -181 1467 -147
rect 1535 -181 1547 -147
rect 1455 -187 1547 -181
rect 1613 -147 1705 -141
rect 1613 -181 1625 -147
rect 1693 -181 1705 -147
rect 1613 -187 1705 -181
rect 1771 -147 1863 -141
rect 1771 -181 1783 -147
rect 1851 -181 1863 -147
rect 1771 -187 1863 -181
rect 1929 -147 2021 -141
rect 1929 -181 1941 -147
rect 2009 -181 2021 -147
rect 1929 -187 2021 -181
rect 2087 -147 2179 -141
rect 2087 -181 2099 -147
rect 2167 -181 2179 -147
rect 2087 -187 2179 -181
rect 2245 -147 2337 -141
rect 2245 -181 2257 -147
rect 2325 -181 2337 -147
rect 2245 -187 2337 -181
rect 2403 -147 2495 -141
rect 2403 -181 2415 -147
rect 2483 -181 2495 -147
rect 2403 -187 2495 -181
rect 2561 -147 2653 -141
rect 2561 -181 2573 -147
rect 2641 -181 2653 -147
rect 2561 -187 2653 -181
rect 2719 -147 2811 -141
rect 2719 -181 2731 -147
rect 2799 -181 2811 -147
rect 2719 -187 2811 -181
rect 2877 -147 2969 -141
rect 2877 -181 2889 -147
rect 2957 -181 2969 -147
rect 2877 -187 2969 -181
rect 3035 -147 3127 -141
rect 3035 -181 3047 -147
rect 3115 -181 3127 -147
rect 3035 -187 3127 -181
rect 3193 -147 3285 -141
rect 3193 -181 3205 -147
rect 3273 -181 3285 -147
rect 3193 -187 3285 -181
rect 3351 -147 3443 -141
rect 3351 -181 3363 -147
rect 3431 -181 3443 -147
rect 3351 -187 3443 -181
rect 3509 -147 3601 -141
rect 3509 -181 3521 -147
rect 3589 -181 3601 -147
rect 3509 -187 3601 -181
rect 3667 -147 3759 -141
rect 3667 -181 3679 -147
rect 3747 -181 3759 -147
rect 3667 -187 3759 -181
rect 3825 -147 3917 -141
rect 3825 -181 3837 -147
rect 3905 -181 3917 -147
rect 3825 -187 3917 -181
rect 3983 -147 4075 -141
rect 3983 -181 3995 -147
rect 4063 -181 4075 -147
rect 3983 -187 4075 -181
rect 4141 -147 4233 -141
rect 4141 -181 4153 -147
rect 4221 -181 4233 -147
rect 4141 -187 4233 -181
rect 4299 -147 4391 -141
rect 4299 -181 4311 -147
rect 4379 -181 4391 -147
rect 4299 -187 4391 -181
rect 4457 -147 4549 -141
rect 4457 -181 4469 -147
rect 4537 -181 4549 -147
rect 4457 -187 4549 -181
rect 4615 -147 4707 -141
rect 4615 -181 4627 -147
rect 4695 -181 4707 -147
rect 4615 -187 4707 -181
rect 4773 -147 4865 -141
rect 4773 -181 4785 -147
rect 4853 -181 4865 -147
rect 4773 -187 4865 -181
rect 4931 -147 5023 -141
rect 4931 -181 4943 -147
rect 5011 -181 5023 -147
rect 4931 -187 5023 -181
rect 5089 -147 5181 -141
rect 5089 -181 5101 -147
rect 5169 -181 5181 -147
rect 5089 -187 5181 -181
rect 5247 -147 5339 -141
rect 5247 -181 5259 -147
rect 5327 -181 5339 -147
rect 5247 -187 5339 -181
rect 5405 -147 5497 -141
rect 5405 -181 5417 -147
rect 5485 -181 5497 -147
rect 5405 -187 5497 -181
rect 5563 -147 5655 -141
rect 5563 -181 5575 -147
rect 5643 -181 5655 -147
rect 5563 -187 5655 -181
rect 5721 -147 5813 -141
rect 5721 -181 5733 -147
rect 5801 -181 5813 -147
rect 5721 -187 5813 -181
rect 5879 -147 5971 -141
rect 5879 -181 5891 -147
rect 5959 -181 5971 -147
rect 5879 -187 5971 -181
rect 6037 -147 6129 -141
rect 6037 -181 6049 -147
rect 6117 -181 6129 -147
rect 6037 -187 6129 -181
rect 6195 -147 6287 -141
rect 6195 -181 6207 -147
rect 6275 -181 6287 -147
rect 6195 -187 6287 -181
rect 6353 -147 6445 -141
rect 6353 -181 6365 -147
rect 6433 -181 6445 -147
rect 6353 -187 6445 -181
rect 6511 -147 6603 -141
rect 6511 -181 6523 -147
rect 6591 -181 6603 -147
rect 6511 -187 6603 -181
rect 6669 -147 6761 -141
rect 6669 -181 6681 -147
rect 6749 -181 6761 -147
rect 6669 -187 6761 -181
rect 6827 -147 6919 -141
rect 6827 -181 6839 -147
rect 6907 -181 6919 -147
rect 6827 -187 6919 -181
rect 6985 -147 7077 -141
rect 6985 -181 6997 -147
rect 7065 -181 7077 -147
rect 6985 -187 7077 -181
rect 7143 -147 7235 -141
rect 7143 -181 7155 -147
rect 7223 -181 7235 -147
rect 7143 -187 7235 -181
rect 7301 -147 7393 -141
rect 7301 -181 7313 -147
rect 7381 -181 7393 -147
rect 7301 -187 7393 -181
rect 7459 -147 7551 -141
rect 7459 -181 7471 -147
rect 7539 -181 7551 -147
rect 7459 -187 7551 -181
rect 7617 -147 7709 -141
rect 7617 -181 7629 -147
rect 7697 -181 7709 -147
rect 7617 -187 7709 -181
rect 7775 -147 7867 -141
rect 7775 -181 7787 -147
rect 7855 -181 7867 -147
rect 7775 -187 7867 -181
rect 7933 -147 8025 -141
rect 7933 -181 7945 -147
rect 8013 -181 8025 -147
rect 7933 -187 8025 -181
rect 8091 -147 8183 -141
rect 8091 -181 8103 -147
rect 8171 -181 8183 -147
rect 8091 -187 8183 -181
rect 8249 -147 8341 -141
rect 8249 -181 8261 -147
rect 8329 -181 8341 -147
rect 8249 -187 8341 -181
rect 8407 -147 8499 -141
rect 8407 -181 8419 -147
rect 8487 -181 8499 -147
rect 8407 -187 8499 -181
rect 8565 -147 8657 -141
rect 8565 -181 8577 -147
rect 8645 -181 8657 -147
rect 8565 -187 8657 -181
rect 8723 -147 8815 -141
rect 8723 -181 8735 -147
rect 8803 -181 8815 -147
rect 8723 -187 8815 -181
rect 8881 -147 8973 -141
rect 8881 -181 8893 -147
rect 8961 -181 8973 -147
rect 8881 -187 8973 -181
rect 9039 -147 9131 -141
rect 9039 -181 9051 -147
rect 9119 -181 9131 -147
rect 9039 -187 9131 -181
rect 9197 -147 9289 -141
rect 9197 -181 9209 -147
rect 9277 -181 9289 -147
rect 9197 -187 9289 -181
rect 9355 -147 9447 -141
rect 9355 -181 9367 -147
rect 9435 -181 9447 -147
rect 9355 -187 9447 -181
rect 9513 -147 9605 -141
rect 9513 -181 9525 -147
rect 9593 -181 9605 -147
rect 9513 -187 9605 -181
rect 9671 -147 9763 -141
rect 9671 -181 9683 -147
rect 9751 -181 9763 -147
rect 9671 -187 9763 -181
rect 9829 -147 9921 -141
rect 9829 -181 9841 -147
rect 9909 -181 9921 -147
rect 9829 -187 9921 -181
rect 9987 -147 10079 -141
rect 9987 -181 9999 -147
rect 10067 -181 10079 -147
rect 9987 -187 10079 -181
rect 10145 -147 10237 -141
rect 10145 -181 10157 -147
rect 10225 -181 10237 -147
rect 10145 -187 10237 -181
rect 10303 -147 10395 -141
rect 10303 -181 10315 -147
rect 10383 -181 10395 -147
rect 10303 -187 10395 -181
rect 10461 -147 10553 -141
rect 10461 -181 10473 -147
rect 10541 -181 10553 -147
rect 10461 -187 10553 -181
rect 10619 -147 10711 -141
rect 10619 -181 10631 -147
rect 10699 -181 10711 -147
rect 10619 -187 10711 -181
rect 10777 -147 10869 -141
rect 10777 -181 10789 -147
rect 10857 -181 10869 -147
rect 10777 -187 10869 -181
rect 10935 -147 11027 -141
rect 10935 -181 10947 -147
rect 11015 -181 11027 -147
rect 10935 -187 11027 -181
rect 11093 -147 11185 -141
rect 11093 -181 11105 -147
rect 11173 -181 11185 -147
rect 11093 -187 11185 -181
rect 11251 -147 11343 -141
rect 11251 -181 11263 -147
rect 11331 -181 11343 -147
rect 11251 -187 11343 -181
rect 11409 -147 11501 -141
rect 11409 -181 11421 -147
rect 11489 -181 11501 -147
rect 11409 -187 11501 -181
rect 11567 -147 11659 -141
rect 11567 -181 11579 -147
rect 11647 -181 11659 -147
rect 11567 -187 11659 -181
rect 11725 -147 11817 -141
rect 11725 -181 11737 -147
rect 11805 -181 11817 -147
rect 11725 -187 11817 -181
rect 11883 -147 11975 -141
rect 11883 -181 11895 -147
rect 11963 -181 11975 -147
rect 11883 -187 11975 -181
rect 12041 -147 12133 -141
rect 12041 -181 12053 -147
rect 12121 -181 12133 -147
rect 12041 -187 12133 -181
rect 12199 -147 12291 -141
rect 12199 -181 12211 -147
rect 12279 -181 12291 -147
rect 12199 -187 12291 -181
rect 12357 -147 12449 -141
rect 12357 -181 12369 -147
rect 12437 -181 12449 -147
rect 12357 -187 12449 -181
rect 12515 -147 12607 -141
rect 12515 -181 12527 -147
rect 12595 -181 12607 -147
rect 12515 -187 12607 -181
rect 12673 -147 12765 -141
rect 12673 -181 12685 -147
rect 12753 -181 12765 -147
rect 12673 -187 12765 -181
rect 12831 -147 12923 -141
rect 12831 -181 12843 -147
rect 12911 -181 12923 -147
rect 12831 -187 12923 -181
rect 12989 -147 13081 -141
rect 12989 -181 13001 -147
rect 13069 -181 13081 -147
rect 12989 -187 13081 -181
rect 13147 -147 13239 -141
rect 13147 -181 13159 -147
rect 13227 -181 13239 -147
rect 13147 -187 13239 -181
rect 13305 -147 13397 -141
rect 13305 -181 13317 -147
rect 13385 -181 13397 -147
rect 13305 -187 13397 -181
rect 13463 -147 13555 -141
rect 13463 -181 13475 -147
rect 13543 -181 13555 -147
rect 13463 -187 13555 -181
rect 13621 -147 13713 -141
rect 13621 -181 13633 -147
rect 13701 -181 13713 -147
rect 13621 -187 13713 -181
rect 13779 -147 13871 -141
rect 13779 -181 13791 -147
rect 13859 -181 13871 -147
rect 13779 -187 13871 -181
rect 13937 -147 14029 -141
rect 13937 -181 13949 -147
rect 14017 -181 14029 -147
rect 13937 -187 14029 -181
rect 14095 -147 14187 -141
rect 14095 -181 14107 -147
rect 14175 -181 14187 -147
rect 14095 -187 14187 -181
rect 14253 -147 14345 -141
rect 14253 -181 14265 -147
rect 14333 -181 14345 -147
rect 14253 -187 14345 -181
rect 14411 -147 14503 -141
rect 14411 -181 14423 -147
rect 14491 -181 14503 -147
rect 14411 -187 14503 -181
rect 14569 -147 14661 -141
rect 14569 -181 14581 -147
rect 14649 -181 14661 -147
rect 14569 -187 14661 -181
rect 14727 -147 14819 -141
rect 14727 -181 14739 -147
rect 14807 -181 14819 -147
rect 14727 -187 14819 -181
rect 14885 -147 14977 -141
rect 14885 -181 14897 -147
rect 14965 -181 14977 -147
rect 14885 -187 14977 -181
rect 15043 -147 15135 -141
rect 15043 -181 15055 -147
rect 15123 -181 15135 -147
rect 15043 -187 15135 -181
rect 15201 -147 15293 -141
rect 15201 -181 15213 -147
rect 15281 -181 15293 -147
rect 15201 -187 15293 -181
rect 15359 -147 15451 -141
rect 15359 -181 15371 -147
rect 15439 -181 15451 -147
rect 15359 -187 15451 -181
rect 15517 -147 15609 -141
rect 15517 -181 15529 -147
rect 15597 -181 15609 -147
rect 15517 -187 15609 -181
rect 15675 -147 15767 -141
rect 15675 -181 15687 -147
rect 15755 -181 15767 -147
rect 15675 -187 15767 -181
<< properties >>
string FIXED_BBOX -15934 -302 15934 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 200 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
